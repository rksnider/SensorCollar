-- RTC_Set.vhd

-- Generated using ACDS version 15.0 145

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity RTC_Set is
	port (
		source_clk : in  std_logic                     := '0'; -- source_clk.clk
		source     : out std_logic_vector(32 downto 0)         --    sources.source
	);
end entity RTC_Set;

architecture rtl of RTC_Set is
	component altsource_probe is
		generic (
			sld_auto_instance_index : string  := "YES";
			sld_instance_index      : integer := 0;
			instance_id             : string  := "NONE";
			probe_width             : integer := 1;
			source_width            : integer := 1;
			source_initial_value    : string  := "0";
			enable_metastability    : string  := "NO"
		);
		port (
			source     : out std_logic_vector(32 downto 0);        -- source
			source_clk : in  std_logic                     := 'X'; -- clk
			source_ena : in  std_logic                     := 'X'  -- source_ena
		);
	end component altsource_probe;

begin

	in_system_sources_probes_0 : component altsource_probe
		generic map (
			sld_auto_instance_index => "NO",
			sld_instance_index      => 0,
			instance_id             => "RTC",
			probe_width             => 0,
			source_width            => 33,
			source_initial_value    => "0",
			enable_metastability    => "YES"
		)
		port map (
			source     => source,     --    sources.source
			source_clk => source_clk, -- source_clk.clk
			source_ena => '1'         -- (terminated)
		);

end architecture rtl; -- of RTC_Set
