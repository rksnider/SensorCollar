----------------------------------------------------------------------------
--
--! @file       Collar.vhd
--! @brief      Acoustic Recording Collar Top Level.
--! @details    Instanciates and connects all the components that make up
--!             the Acoustic Recording Collar FPGA implementation.
--! @author     Emery Newlon
--! @date       March 2015
--! @copyright  Copyright (C) 2015 Ross K. Snider and Emery L. Newlon
--
--  This program is free software: you can redistribute it and/or modify
--  it under the terms of the GNU General Public License as published by
--  the Free Software Foundation, either version 3 of the License, or
--  (at your option) any later version.
--
--  This program is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--  GNU General Public License for more details.
--
--  You should have received a copy of the GNU General Public License
--  along with this program.  If not, see <http://www.gnu.org/licenses/>.
--
--  Emery Newlon
--  Electrical and Computer Engineering
--  Montana State University
--  610 Cobleigh Hall
--  Bozeman, MT 59717
--  emery.newlon@msu.montana.edu
--
----------------------------------------------------------------------------

library IEEE ;                  --! Use standard library.
use IEEE.STD_LOGIC_1164.ALL ;   --! Use standard logic elements.
use IEEE.NUMERIC_STD.ALL ;      --! Use numeric standard.
use IEEE.MATH_REAL.ALL ;        --! Real number functions.

library GENERAL ;               --! General libraries
use GENERAL.UTILITIES_PKG.ALL ;

library WORK ;                  --! Local libraries
use WORK.PC_STATUSCONTROL_PKG.ALL ;
use WORK.SDRAM_INFORMATION_PKG.ALL ;


----------------------------------------------------------------------------
--
--! @brief      Acoustic Recording Collar Top Level.
--! @details    Instanciates and connects all the components that make up
--!             the Acoustic Recording Collar FPGA implementation.
--!
--! @param      master_clk_freq_g Frequency of the system clock in cycles
--!                               per second.
--! @param      button_cnt_g    Number of buttons used by the device.
--! @param      master_clk      Clock generated by the system that drives
--!                             everything else.
--! @param      buttons_in      Vector of button signals used by the device.
--! @param      sdram_clk         Clock driving the SDRAM.
--! @param      sdram_clk_en_out  The clock is enabled on the SDRAM.
--! @param      sdram_command_out The command sent to the SDRAM.
--! @param      sdram_mask_out    The bytes masked from the SDRAM data bus.
--! @param      sdram_bank_out    The SDRAM bank to access.
--! @param      sdram_addr_out    The SDRAM row or column to access.
--! @param      sdram_data_io     The SDRAM data bus.
--! @param      log_*             These pins miror the other pins for
--!                               logging to test points.
--! @param      log_empty_out     The SDRAM and buffers are empty.
--! @param      log_forceout_out  Forcing output of the SDRAM.
--! @param      log_fail_out      The input from SDRAM did not match the
--!                               expected input.
--
----------------------------------------------------------------------------

entity SDRAM_ControllerTest_tb is

  Generic (
    master_clk_freq_g     : natural   := 10e6 ;
    button_cnt_g          : natural   :=  8
  ) ;
  Port (
    master_clk            : in    std_logic ;
    buttons_in            : in    std_logic_vector (button_cnt_g-1
                                                    downto 0) ;

    sdram_clk             : out   std_logic ;
    sdram_clk_en_out      : out   std_logic ;
    sdram_command_out     : out   std_logic_vector (3 downto 0) ;
    sdram_mask_out        : out   std_logic_vector (1 downto 0) ;
    sdram_bank_out        : out   std_logic_vector (1 downto 0) ;

    sdram_addr_out        : out   std_logic_vector (12 downto 0) ;
    sdram_data_io         : inout std_logic_vector (15 downto 0) ;

    PC_StatusChg_in       : in    std_logic ;
    PC_SPI_clk_out        : out   std_logic ;
    PC_SPI_mosi_out       : out   std_logic ;
    PC_SPI_miso_in        : in    std_logic ;
    PC_SPI_cs_n_out       : out   std_logic ;

    log_clk_out           : out   std_logic ;
    log_clk_en_out        : out   std_logic ;
    log_command_out       : out   std_logic_vector (3 downto 0) ;
    log_mask_out          : out   std_logic_vector (1 downto 0) ;
    log_bank_out          : out   std_logic_vector (1 downto 0) ;
    log_addr_out          : out   std_logic_vector (12 downto 0) ;
    log_data_out          : out   std_logic_vector (15 downto 0) ;
    log_empty_out         : out   std_logic ;
    log_forceout_out      : out   std_logic ;
    log_fail_out          : out   std_logic

  ) ;

end entity SDRAM_ControllerTest_tb ;


architecture rtl of SDRAM_ControllerTest_tb is

  --  Memory components.

  constant outmem_bytecnt_c     : natural := 4096 ;
  constant outmem_rdwidth_c     : natural := 32 ;
  constant outmem_wrwidth_c     : natural := 16 ;
  constant outmem_buffcount_c   : natural := 2 ;

  constant outmem_rdaddrbits_c  : natural :=
              const_bits ((8 * outmem_bytecnt_c / outmem_rdwidth_c) - 1) ;
  constant outmem_wraddrbits_c  : natural :=
              const_bits ((8 * outmem_bytecnt_c / outmem_wrwidth_c) - 1) ;

  component outmem IS
    PORT
    (
      data        : IN STD_LOGIC_VECTOR (outmem_wrwidth_c-1 DOWNTO 0) ;
      rdaddress   : IN STD_LOGIC_VECTOR (outmem_rdaddrbits_c-1 DOWNTO 0) ;
      rdclock     : IN STD_LOGIC ;
      rden        : IN STD_LOGIC  := '1' ;
      wraddress   : IN STD_LOGIC_VECTOR (outmem_wraddrbits_c-1 DOWNTO 0) ;
      wrclock     : IN STD_LOGIC  := '1' ;
      wren        : IN STD_LOGIC  := '0' ;
      q           : OUT STD_LOGIC_VECTOR (outmem_rdwidth_c-1 DOWNTO 0)
    ) ;
  END component outmem ;

  constant inmem_bytecnt_c      : natural := 4096 ;
  constant inmem_rdwidth_c      : natural := 16 ;
  constant inmem_wrwidth_c      : natural := 32 ;
  constant inmem_buffcount_c    : natural := 2 ;

  constant inmem_rdaddrbits_c   : natural :=
              const_bits ((8 * inmem_bytecnt_c / inmem_rdwidth_c) - 1) ;
  constant inmem_wraddrbits_c   : natural :=
              const_bits ((8 * inmem_bytecnt_c / inmem_wrwidth_c) - 1) ;

  component inmem IS
    PORT
    (
      data        : IN STD_LOGIC_VECTOR (inmem_wrwidth_c-1 DOWNTO 0) ;
      rdaddress   : IN STD_LOGIC_VECTOR (inmem_rdaddrbits_c-1 DOWNTO 0) ;
      rdclock     : IN STD_LOGIC ;
      rden        : IN STD_LOGIC  := '1' ;
      wraddress   : IN STD_LOGIC_VECTOR (inmem_wraddrbits_c-1 DOWNTO 0) ;
      wrclock     : IN STD_LOGIC  := '1' ;
      wren        : IN STD_LOGIC  := '0' ;
      q           : OUT STD_LOGIC_VECTOR (inmem_rdwidth_c-1 DOWNTO 0)
    ) ;
  END component inmem ;

  --  SDRAM controller componenent.

  component SDRAM_Controller is

    Generic (
      sysclk_freq_g         : natural     := 10e6 ;

      outmem_buffrows_g     : natural     := 1 ;
      outmem_buffcount_g    : natural     := 2 ;
      inmem_buffouts_g      : natural     := 1 ;
      inmem_buffcount_g     : natural     := 2 ;
      sdram_space_g         : SDRAM_Capacity_t  := SDRAM_32_Capacity_c ;
      sdram_times_g         : SDRAM_Timing_t    := SDRAM_75_3_Timing_c
    ) ;
    Port (
      reset                 : in    std_logic ;
      sysclk                : in    std_logic ;

      ready_out             : out   std_logic ;

      inmem_buffready_in    : in    std_logic ;
      inmem_datafrom_in     : in    std_logic_vector (sdram_space_g.DATABITS-1
                                                      downto 0) ;
      inmem_address_out     : out
          std_logic_vector (const_bits (inmem_buffcount_g * inmem_buffouts_g *
                                        outmem_buffrows_g *
                                        sdram_space_g.ROWBITS /
                                        sdram_space_g.DATABITS - 1) - 1
                                          downto 0) ;
      inmem_read_en_out     : out   std_logic ;
      inmem_clk_out         : out   std_logic ;

      outmem_buffready_in   : in    std_logic ;
      outmem_datato_out     : out   std_logic_vector (sdram_space_g.DATABITS-1
                                                      downto 0) ;
      outmem_address_out    : out
          std_logic_vector (const_bits (outmem_buffcount_g *
                                        outmem_buffrows_g *
                                        sdram_space_g.ROWBITS /
                                        sdram_space_g.DATABITS - 1) - 1
                                          downto 0) ;
      outmem_write_en_out   : out   std_logic ;
      outmem_clk_out        : out   std_logic ;
      outmem_amt_out        : out
          unsigned (const_bits (sdram_space_g.BANKS * sdram_space_g.ROWCOUNT *
                                sdram_space_g.ROWBITS / 8 - 1) - 1 downto 0) ;
      outmem_writing_out    : out   std_logic ;

      sdram_data_in         : in    std_logic_vector (sdram_space_g.DATABITS-1
                                                        downto 0) ;
      sdram_data_out        : out   std_logic_vector (sdram_space_g.DATABITS-1
                                                        downto 0) ;
      sdram_data_dir        : out   std_logic ;

      sdram_mask_out        : out
          std_logic_vector (sdram_space_g.DATABITS / 8 - 1 downto 0) ;
      sdram_address_out     : out   unsigned (sdram_space_g.ADDRBITS-1
                                                        downto 0) ;
      sdram_bank_out        : out
          unsigned (const_bits (sdram_space_g.BANKS - 1)-1 downto 0) ;
      sdram_command_out     : out   std_logic_vector (sdram_space_g.CMDBITS-1
                                                        downto 0) ;
      sdram_clk_en_out      : out   std_logic ;
      sdram_clk_out         : out   std_logic ;
      sdram_empty_out       : out   std_logic ;
      sdram_forceout_in     : in    std_logic
    ) ;

  end component SDRAM_Controller ;

  --  Global nternal clock.

  constant clk_freq_target_c  : natural := 1e6 ;

  constant clk_count_c        : natural :=
        natural (trunc (real (master_clk_freq_g) /
                        real (clk_freq_target_c) / 2.0 + 0.5)) ;

  constant clk_freq_c         : natural :=
        natural (trunc (real (master_clk_freq_g) /
                        real (clk_count_c) / 2.0)) ;

  signal int_clk_count        : unsigned (const_bits (clk_count_c-1) - 1
                                          downto 0) ;

  signal internal_clk         : std_logic ;
  signal global_int_clk       : std_logic ;

  -- attribute keep                    : boolean ;
  -- attribute keep of global_int_clk  : signal is true ;

  component internal_clock is
  port (
    inclk            : IN    STD_LOGIC ;
    outclk           : OUT   STD_LOGIC
  ) ;
  end component internal_clock ;

  --  Power Controller SPI communications channel.

  constant cs_sdram_set_c         : ControlSignalsArray :=
  (
    Ctl_SDRAM_On_e,
    Ctl_SDRAM_On_e
  ) ;

  signal PC_StatusReg             : std_logic_vector (StatusSignalsCnt_c-1
                                                      downto 0) ;
  signal PC_StatusSet             : std_logic ;
  signal PC_ControlReg            : std_logic_vector (ControlSignalsCnt_c-1
                                                      downto 0) :=
                                        controlSignalsSet (cs_sdram_set_c) ;

  component StatCtlSPI_FPGA is
    Generic (
      status_bits_g               : natural := 16 ;
      control_bits_g              : natural := 16 ;
      flash_bytes_transfer        : natural := 0 ;
      data_length_bit_width_g     : natural := 8
    ) ;
    Port (
      clk                         : in    std_logic ;
      rst_n                       : in    std_logic ;
      status_out                  : out   std_logic_vector (status_bits_g-1
                                                            downto 0) ;
      status_chg_in               : in    std_logic ;
      status_set_out              : out   std_logic ;
      control_in                  : in    std_logic_vector (control_bits_g-1
                                                            downto 0) ;

      sclk                        : out   std_logic ;
      mosi                        : out   std_logic ;
      miso                        : in    std_logic ;
      cs_n                        : out   std_logic
    ) ;
  end component StatCtlSPI_FPGA ;

  --  Button specifications.

  constant reset_button_c   : natural := 0 ;

  --  Reset information.  The power up signal defaults to zero.

  constant pu_count_c       : natural := 3 ;

  signal reset              : std_logic ;
  signal power_up           : std_logic := '0' ;
  signal pu_counter         : unsigned (const_bits (pu_count_c)-1
                                        downto 0) := (others => '0') ;

  constant pb_time_c        : real    := 0.5 ;
  constant pb_count_c       : natural :=
              natural (trunc (real (master_clk_freq_g) * pb_time_c)) ;
  constant pb_count_bits_c  : natural := const_bits (pb_count_c) ;

  signal reset_pushed       : std_logic := '0' ;
  signal pb_counter         : unsigned (pb_count_bits_c-1 downto 0) :=
                                (others => '0') ;

  --  SDRAM information.

  constant sdram_space_c        : SDRAM_Capacity_t := SDRAM_16_Capacity_c ;

  --  Buffer dual port RAM communication signals.

  constant outmem_buffbytes_c     : natural :=
              (outmem_bytecnt_c / outmem_buffcount_c) ;
  constant outmem_buffrows_c      : natural :=
              (outmem_buffbytes_c / (sdram_space_c.ROWBITS / 8)) ;

  signal outmem_read_addr         : std_logic_vector (outmem_rdaddrbits_c-1
                                                      downto 0) ;
  signal outmem_read_clk          : std_logic ;
  signal outmem_read_en           : std_logic ;
  signal outmem_read_data         : std_logic_vector (outmem_rdwidth_c-1
                                                      downto 0) ;

  signal outmem_write_addr        : std_logic_vector (outmem_wraddrbits_c-1
                                                      downto 0) ;
  signal outmem_write_clk         : std_logic ;
  signal outmem_write_en          : std_logic ;
  signal outmem_write_data        : std_logic_vector (outmem_wrwidth_c-1
                                                      downto 0) ;

  signal outmem_write_amt         :
            unsigned (const_bits (sdram_space_c.BANKS *
                                  sdram_space_c.ROWCOUNT *
                                  sdram_space_c.ROWBITS / 8 - 1) - 1
                      downto 0) ;
  signal outmem_writing           : std_logic ;
  signal outmem_writing_fwl       : std_logic ;
  signal outmem_buff_ready        : std_logic ;

  signal reading_amt              : unsigned (outmem_write_amt'length-1
                                              downto 0) ;
  signal reading_done             : unsigned (reading_amt'length-1
                                              downto 0) ;
  signal reading_active           : std_logic ;

  constant outmem_interval_c      : natural :=
              natural (0.001 * real (clk_freq_c)) ;

  signal outmem_timer             :
              unsigned (const_bits (outmem_interval_c) - 1 downto 0) ;
  signal output_count             : unsigned (31 downto 0) ;

  signal output_fail_read         : unsigned (31 downto 0) ;
  signal output_fail_cnt          : unsigned (31 downto 0) ;

  constant inmem_buffbytes_c      : natural :=
              (inmem_bytecnt_c / inmem_buffcount_c) ;
  constant inmem_buffouts_c       : natural :=
              (outmem_buffbytes_c / inmem_buffbytes_c) ;

  signal inmem_read_addr          : std_logic_vector (inmem_rdaddrbits_c-1
                                                      downto 0) ;
  signal inmem_read_clk           : std_logic ;
  signal inmem_read_en            : std_logic ;
  signal inmem_read_data          : std_logic_vector (inmem_rdwidth_c-1
                                                      downto 0) ;

  signal inmem_write_addr         : std_logic_vector (inmem_wraddrbits_c-1
                                                      downto 0) ;
  signal inmem_write_clk          : std_logic ;
  signal inmem_write_en           : std_logic ;
  signal inmem_write_data         : std_logic_vector (inmem_wrwidth_c-1
                                                      downto 0) ;

  constant inmem_interval_c       : natural :=
              natural (0.030 * real (clk_freq_c)) ;

  signal inmem_count              : unsigned (31 downto 0) ;
  signal inmem_timer              :
            unsigned (const_bits (inmem_interval_c) - 1 downto 0) ;
  signal inmem_buff_ready         : std_logic ;

  --  SDRAM signals.

  signal sdram_data_from      : std_logic_vector (sdram_space_c.DATABITS-1
                                                  downto 0) ;
  signal sdram_data_to        : std_logic_vector (sdram_space_c.DATABITS-1
                                                  downto 0) ;
  signal sdram_data_drive     : std_logic ;
  signal sdram_mask           :
            std_logic_vector (sdram_space_c.DATABITS / 8 - 1 downto 0) ;
  signal sdram_address        : unsigned (sdram_space_c.ADDRBITS-1
                                          downto 0) ;
  signal sdram_bank           :
            unsigned (const_bits (sdram_space_c.BANKS-1) - 1 downto 0) ;
  signal sdram_command        : std_logic_vector (sdram_space_c.CMDBITS-1
                                                  downto 0) ;
  signal sdram_clk_en         : std_logic ;
  signal sdram_clock          : std_logic ;
  signal sdram_empty          : std_logic ;
  signal sdram_forceout       : std_logic ;
  signal sdram_ready          : std_logic ;


begin

  --------------------------------------------------------------------------
  --  Memory instances.
  --------------------------------------------------------------------------

  input_mem : inmem
    port map
    (
      rdaddress   => inmem_read_addr,
      rdclock     => inmem_read_clk,
      rden        => inmem_read_en,
      q           => inmem_read_data,
      wraddress   => inmem_write_addr,
      wrclock     => inmem_write_clk,
      wren        => inmem_write_en,
      data        => inmem_write_data
    ) ;

  output_mem : outmem
    port map
    (
      rdaddress   => outmem_read_addr,
      rdclock     => outmem_read_clk,
      rden        => outmem_read_en,
      q           => outmem_read_data,
      wraddress   => outmem_write_addr,
      wrclock     => outmem_write_clk,
      wren        => outmem_write_en,
      data        => outmem_write_data
    ) ;

  outmem_read_en            <= '1' ;

  --------------------------------------------------------------------------
  --  Power Controller SPI communications channel instance.
  --------------------------------------------------------------------------

  pc_spi : StatCtlSPI_FPGA
    Generic Map (
      status_bits_g               => StatusSignalsCnt_c,
      control_bits_g              => ControlSignalsCnt_c,
      flash_bytes_transfer        => 0,
      data_length_bit_width_g     => 8
    )
    Port Map (
      clk                         => global_int_clk,
      rst_n                       => not reset,
      status_out                  => PC_StatusReg,
      status_chg_in               => PC_StatusChg_in,
      status_set_out              => PC_StatusSet,
      control_in                  => PC_ControlReg,

      sclk                        => PC_SPI_clk_out,
      mosi                        => PC_SPI_mosi_out,
      miso                        => PC_SPI_miso_in,
      cs_n                        => PC_SPI_cs_n_out
    ) ;

  --------------------------------------------------------------------------
  --  SDRAM controller instance.
  --------------------------------------------------------------------------

  sdram_ctl : SDRAM_Controller

    Generic Map (
      sysclk_freq_g         => clk_freq_c,

      outmem_buffrows_g     => outmem_buffrows_c,
      outmem_buffcount_g    => outmem_buffcount_c,
      inmem_buffouts_g      => inmem_buffouts_c,
      inmem_buffcount_g     => inmem_buffcount_c,
      sdram_space_g         => sdram_space_c,
      sdram_times_g         => SDRAM_75_3_Timing_c
    )
    Port Map (
      reset                 => reset,
      sysclk                => global_int_clk,

      ready_out             => sdram_ready,

      inmem_buffready_in    => inmem_buff_ready,
      inmem_datafrom_in     => inmem_read_data,
      inmem_address_out     => inmem_read_addr,
      inmem_read_en_out     => inmem_read_en,
      inmem_clk_out         => inmem_read_clk,

      outmem_buffready_in   => outmem_buff_ready,
      outmem_datato_out     => outmem_write_data,
      outmem_address_out    => outmem_write_addr,
      outmem_write_en_out   => outmem_write_en,
      outmem_clk_out        => outmem_write_clk,
      outmem_amt_out        => outmem_write_amt,
      outmem_writing_out    => outmem_writing,

      sdram_data_in         => sdram_data_from,
      sdram_data_out        => sdram_data_to,
      sdram_data_dir        => sdram_data_drive,

      sdram_mask_out        => sdram_mask,
      sdram_address_out     => sdram_address,
      sdram_bank_out        => sdram_bank,
      sdram_command_out     => sdram_command,
      sdram_clk_en_out      => sdram_clk_en,
      sdram_clk_out         => sdram_clock,
      sdram_empty_out       => sdram_empty,
      sdram_forceout_in     => sdram_forceout
    ) ;

  sdram_data_io       <= sdram_data_to when (sdram_data_drive = '1') else
                         (others => 'Z') ;
  sdram_data_from     <= sdram_data_io ;

  sdram_clk           <= sdram_clock ;
  sdram_clk_en_out    <= sdram_clk_en ;
  sdram_command_out   <= sdram_command ;
  sdram_mask_out      <= sdram_mask ;
  sdram_bank_out      <= std_logic_vector (sdram_bank) ;
  sdram_addr_out      <= std_logic_vector (sdram_address) ;

  log_data_out        <= sdram_data_to ;
  log_clk_out         <= sdram_clock ;
  log_clk_en_out      <= sdram_clk_en ;
  log_command_out     <= sdram_command ;
  log_mask_out        <= sdram_mask ;
  log_bank_out        <= std_logic_vector (sdram_bank) ;
  log_addr_out        <= std_logic_vector (sdram_address) ;
  log_empty_out       <= sdram_empty ;
  log_forceout_out    <= sdram_forceout ;

  sdram_forceout      <= '0' ;

  --------------------------------------------------------------------------
  --  Reset occurs on power up or button press of the reset button.
  --------------------------------------------------------------------------

  reset                     <= (not power_up) or reset_pushed ;

  reset_poweron : process (master_clk)
  begin
    if (rising_edge (master_clk)) then
      if (pu_counter = pu_count_c) then
        power_up              <= '1' ;
      else
        pu_counter            <= pu_counter + 1 ;
      end if ;
    end if ;
  end process reset_poweron ;

  --  Debounce the reset button by making sure it is held up or down for a
  --  long period of time.

  reset_pb : process (master_clk)
  begin
    if (rising_edge (master_clk)) then

      if (buttons_in (reset_button_c) /= reset_pushed) then
        if (pb_counter = pb_count_c) then
          reset_pushed      <= buttons_in (reset_button_c) ;
          pb_counter        <= (others => '0') ;
        else
          pb_counter        <= pb_counter + 1 ;
        end if ;
      else
        pb_counter          <= (others => '0') ;
      end if ;
    end if ;
  end process reset_pb ;

  --------------------------------------------------------------------------
  --  Generate internal clock.
  --------------------------------------------------------------------------

  gbl_intclk : internal_clock
  port map (
    inclk                => internal_clk,
    outclk              => global_int_clk
  ) ;

  gen_clock : process (reset, master_clk)
  begin
    if (reset = '1') then
      internal_clk      <= '0' ;
      int_clk_count     <= (others => '0') ;

    elsif (rising_edge (master_clk)) then
      if (int_clk_count /= clk_count_c - 1) then
        int_clk_count   <= int_clk_count + 1 ;
      else
        int_clk_count   <= (others => '0') ;
        internal_clk    <= not internal_clk ;
      end if ;
    end if ;
  end process gen_clock ;

  --------------------------------------------------------------------------
  --  Periodically write a set of sequencial numbers to an input buffer.
  --------------------------------------------------------------------------

  inmem_write_clk           <= not global_int_clk ;

  inmem_fill : process (reset, global_int_clk)
  begin
    if (reset = '1') then
      inmem_count           <= (others => '0') ;
      inmem_timer           <= (others => '0') ;
      inmem_write_addr      <= (others => '1') ;    --  minus one
      inmem_buff_ready      <= '0' ;

    elsif (rising_edge (global_int_clk)) then
      inmem_write_en        <= '0' ;
      inmem_buff_ready      <= '0' ;

      if (sdram_ready = '1') then
        --  Periodically fill an input buffer.

        if (inmem_timer /= inmem_interval_c) then
          inmem_timer         <= inmem_timer + 1 ;
        else
          if ((unsigned (inmem_write_addr) and
               TO_UNSIGNED (inmem_buffbytes_c - 1,
                            inmem_write_addr'length)) =
              TO_UNSIGNED (inmem_buffbytes_c - 2,
                           inmem_write_addr'length)) then

            inmem_timer       <= (others => '0') ;
            inmem_buff_ready  <= '1' ;
          end if ;

          inmem_write_data  <= std_logic_vector (inmem_count) ;
          inmem_write_addr  <= std_logic_vector (
                                    unsigned (inmem_write_addr) + 1) ;
          inmem_write_en    <= '1' ;
          inmem_count       <= inmem_count + 1 ;
        end if ;
      end if ;
    end if ;
  end process inmem_fill ;

  --------------------------------------------------------------------------
  --  Periodically read a set of sequencials number from an output buffer.
  --------------------------------------------------------------------------

  outmem_read_clk               <= not global_int_clk ;

  outmem_empty : process (reset, global_int_clk)
  begin
    if (reset = '1') then
      output_count              <= (others => '0') ;
      outmem_timer              <= (others => '0') ;
      outmem_read_addr          <= (others => '0') ;
      outmem_buff_ready         <= '0' ;
      outmem_writing_fwl        <= '0' ;
      reading_active            <= '0' ;
      reading_amt               <= (others => '0') ;
      reading_done              <= (others => '0') ;
      log_fail_out              <= '0' ;

    elsif (rising_edge (global_int_clk)) then
      outmem_buff_ready         <= '0' ;

      --  Activate reading when signalled to.

      if (sdram_ready = '1') then
        if (outmem_writing_fwl /= outmem_writing) then
          outmem_writing_fwl      <= outmem_writing ;

          if (outmem_writing = '1') then
            reading_active        <= '1' ;
            reading_amt           <= outmem_write_amt ;
            reading_done          <= (others => '0') ;
          end if ;
        end if ;

        if (reading_active = '1') then
          if (reading_amt = reading_done) then
            reading_active        <= '0' ;

          else
            --  Periodically read an output buffer.

            if (outmem_timer /= outmem_interval_c) then
              outmem_timer        <= outmem_timer + 1 ;
            else
              if ((unsigned (outmem_read_addr) and
                   TO_UNSIGNED (outmem_buffbytes_c - 1,
                                outmem_read_addr'length)) =
                  TO_UNSIGNED (outmem_buffbytes_c - 1,
                               outmem_read_addr'length)) then

                reading_done      <= reading_done + outmem_buffbytes_c ;
                outmem_timer      <= (others => '0') ;
                outmem_buff_ready <= '1' ;
              end if ;

              if (unsigned (outmem_read_data) /= output_count) then
                output_fail_read  <= unsigned (outmem_read_data) ;
                output_fail_cnt   <= output_count ;
                log_fail_out      <= '1' ;
              end if ;

              outmem_read_addr    <= std_logic_vector (
                                          unsigned (outmem_read_addr) + 1) ;
              output_count        <= output_count + 1 ;
            end if ;
          end if ;
        end if ;
      end if ;
    end if ;
  end process outmem_empty ;


end architecture rtl ;
