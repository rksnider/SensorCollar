----------------------------------------------------------------------------
--
--! @file       Collar.vhd
--! @brief      Acoustic Recording Collar Top Level.
--! @details    Instanciates and connects all the components that make up
--!             the Acoustic Recording Collar FPGA implementation.
--! @author     Emery Newlon
--! @date       August 2014
--! @copyright  Copyright (C) 2014 Ross K. Snider and Emery L. Newlon
--
--  This program is free software: you can redistribute it and/or modify
--  it under the terms of the GNU General Public License as published by
--  the Free Software Foundation, either version 3 of the License, or
--  (at your option) any later version.
--
--  This program is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--  GNU General Public License for more details.
--
--  You should have received a copy of the GNU General Public License
--  along with this program.  If not, see <http://www.gnu.org/licenses/>.
--
--  Emery Newlon
--  Electrical and Computer Engineering
--  Montana State University
--  610 Cobleigh Hall
--  Bozeman, MT 59717
--  emery.newlon@msu.montana.edu
--
----------------------------------------------------------------------------

library IEEE ;                  --! Use standard library.
use IEEE.STD_LOGIC_1164.ALL ;   --! Use standard logic elements.
use IEEE.NUMERIC_STD.ALL ;      --! Use numeric standard.
use IEEE.MATH_REAL.ALL ;        --! Real number functions.

LIBRARY lpm ;                   --  Use Library of Parameterized Modules.
USE lpm.lpm_components.all ;

library GENERAL ;               --! General libraries
use GENERAL.UTILITIES_PKG.ALL ;

use GENERAL.GPS_CLOCK_PKG.ALL ;
use GENERAL.FORMATSECONDS_PKG.ALL ;

library WORK ;                  --! Local Library
use WORK.COLLAR_CONTROL_PKG.ALL ;
use WORK.COLLAR_PARAMETERS_PKG.ALL ;
use WORK.COLLAR_EVENTS_PKG.ALL ;
use WORK.SHARED_SDC_VALUES_PKG.ALL ;
use WORK.PC_STATUSCONTROL_PKG.ALL ;
use WORK.SDRAM_INFORMATION_PKG.ALL ;
use WORK.MAGMEM_BUFFER_DEF_PKG.ALL ;

use WORK.GPS_MESSAGE_CTL_PKG.ALL ;
use WORK.MSG_UBX_NAV_SOL_PKG.ALL ;
use WORK.MSG_UBX_TIM_TM2_PKG.ALL ;


----------------------------------------------------------------------------
--
--! @brief      Acoustic Recording Collar Top Level.
--! @details    Instanciates and connects all the components that make up
--!             the Acoustic Recording Collar FPGA implementation.
--!
--! @param      source_clk_freq_g Frequency of the system clock in cycles
--!                               per second.
--! @param      button_cnt_g    Number of buttons used by the device.
--! @param      sdram_space_g   Space available parameters for SDRAM chip.
--! @param      sdram_times_g   Timing limits for SDRAM chip.
--! @param      source_clk      Clock generated by the system that drives
--!                             everything else.
--! @param      buttons_in      Vector of button signals used by the device.
--! @param      batt_int_in     Battery monitor interrupt signal.
--! @param      forced_start_in A forced startup has been initiated.
--! @param      i2c_clk_io      I2C bus clock is input or output depending
--!                             on the device driving it.
--! @param      i2c_data_io     I2C bus data is driven by the same device
--!                             that is driving the clock.
--! @param      pc_statchg_in   The Power Controller status register has
--!                             changed and should be reloaded.
--! @param      pc_spi_clk      The Power Controller status register/
--!                             control register SPI bus clock.
--! @param      pc_spi_cs_out   The PC SPI bus chip select.  An SPI
--!                             transfer is initiated when it goes high.
--! @param      pc_spi_mosi_out Master Out/Slave In SPI data line.
--! @param      pc_spi_miso_in  Master In/Slave Out SPI data line.
--! @param      pc_flash_clk      Power Controller Flash access clock.
--! @param      pc_flash_cs_out   PC Flash chip select.
--! @param      pc_flash_data_io  PC Flash data bus.
--! @param      pc_flash_dir_out  PC Flash data direction.  The PC Flash
--!                               bus is high impedance when this line is
--!                               low, driven when it is high.
--! @param      sdram_clk         Clock driving the SDRAM.
--! @param      sdram_clk_en_out  The clock is enabled on the SDRAM.
--! @param      sdram_command_out The command sent to the SDRAM.
--! @param      sdram_mask_out    The bytes masked from the SDRAM data bus.
--! @param      sdram_bank_out    The SDRAM bank to access.
--! @param      sdram_addr_out    The SDRAM row or column to access.
--! @param      sdram_data_io     The SDRAM data bus.
--! @param      sd_clk          Micro SDCard clock.
--! @param      sd_cmd_io       Command line used with the micro SDCard.
--! @param      sd_data_io      Data lines used with the micro SDCard.
--! @param      sdh_clk         High voltage micro SDCard clock.
--! @param      sdh_cmd_io      High voltage command line used with the
--!                             micro SDCard.
--! @param      sdh_data_io     High voltage data lines used with the micro
--!                             SDCard.
--! @param      gps_rx_io       Receive line from the GPS UART.
--! @param      gps_tx_out      Transmit line to the GPS UART.
--! @param      gps_timemark_out  Time mark generator line to the GPS
--!                               external interrupt.
--! @param      gps_timepulse_io  Time pulse signal from GPS.
--! @param      ms_clk          Motion sensor SPI Clock.
--! @param      ms_mosi_out     Motion sensor SPI Master Out/Slave In.
--! @param      ms_miso_in      Motion sensor SPI Master In/Slave Out.
--! @param      ms_int_in       Motion sensor Interrupt.
--! @param      ms_cs_accgyro_out   Motion sensor A/G SPI chip select.
--! @param      ms_miso_accgyro_io  Motion sensor A/G SPI Master In/Slave
--!                                 Out.
--! @param      ms_int1_accgyro_io  Motion sensor A/G Interrupt 1.
--! @param      ms_int2_accgyro_io  Motion sensor A/G Interrupt 2.
--! @param      ms_cs_mag_out   Motion sensor magnetic SPI chip select.
--! @param      ms_miso_mag_io  Motion sensor magnetic SPI Master In/
--!                             Slave Out.
--! @param      ms_int_mag_io   Motion sensor magnetic Interrupt.
--! @param      ms_drdy_mag_io  Motion sensor magnetic Data Ready.
--! @param      magram_clk            Magnetic RAM SPI clock.
--! @param      magram_cs_out         Magnetic RAM chip select.
--! @param      magram_mosi_out       Magnetic RAM SPI Master Out/Slave In.
--! @param      magram_miso_io        Magnetic RAM SPI Master In/Slave Out.
--! @param      magram_writeprot_out  Magnetic RAM write protect.
--! @param      mic_clk         Microphone clock.
--! @param      mic_right_io    Right microphone data.
--! @param      mic_left_io     Left microphone data.
--! @param      radio_clk       Radio trx/rcv bus clock.
--! @param      radio_data_io   Radio data bus.
--
----------------------------------------------------------------------------

entity Collar is

  Generic (
    source_clk_freq_g     : natural           := 10e6 ;
    button_cnt_g          : natural           :=  8 ;
    sdram_space_g         : SDRAM_Capacity_t  := SDRAM_16_Capacity_c ;
    sdram_times_g         : SDRAM_Timing_t    := SDRAM_75_2_Timing_c
  ) ;
  Port (
    source_clk            : in    std_logic ;
    buttons_in            : in    std_logic_vector (button_cnt_g-1
                                                      downto 0) ;

    batt_int_in           : in    std_logic ;
    forced_start_in       : in    std_logic ;

    i2c_clk_io            : inout std_logic ;
    i2c_data_io           : inout std_logic ;

    pc_statchg_in         : in    std_logic ;
    pc_spi_clk            : out   std_logic ;
    pc_spi_cs_out         : out   std_logic ;
    pc_spi_mosi_out       : out   std_logic ;
    pc_spi_miso_in        : in    std_logic ;

    pc_flash_clk          : out   std_logic ;
    pc_flash_cs_out       : out   std_logic ;
    pc_flash_data_io      : inout std_logic_vector (3 downto 0) ;
    pc_flash_dir_out      : out   std_logic ;

    sdram_clk             : out   std_logic ;
    sdram_clk_en_out      : out   std_logic ;
    sdram_command_out     : out   std_logic_vector (3 downto 0) ;
    sdram_mask_out        : out   std_logic_vector (1 downto 0) ;
    sdram_bank_out        : out   std_logic_vector (1 downto 0) ;

    sdram_addr_out        : out   std_logic_vector (12 downto 0) ;
    sdram_data_io         : inout std_logic_vector (15 downto 0) ;

    sd_clk                : out   std_logic ;
    sd_cmd_io             : inout std_logic ;
    sd_data_io            : inout std_logic_vector (3 downto 0) ;

    sdh_clk               : out   std_logic ;
    sdh_cmd_io            : inout std_logic ;
    sdh_data_io           : inout std_logic_vector (3 downto 0) ;

    gps_rx_io             : inout std_logic ;
    gps_tx_out            : out   std_logic ;
    gps_timemark_out      : out   std_logic ;
    gps_timepulse_io      : inout std_logic ;

    ms_clk                : out   std_logic ;
    ms_mosi_out           : out   std_logic ;
    --ms_miso_in            : in    std_logic ;
    --ms_int_in             : in    std_logic ;

    ms_cs_accgyro_out     : out   std_logic ;
    ms_miso_accgyro_io    : inout std_logic ;
    ms_int1_accgyro_io    : inout std_logic ;
    ms_int2_accgyro_io    : inout std_logic ;

    ms_cs_mag_out         : out   std_logic ;
    ms_miso_mag_io        : inout std_logic ;
    ms_int_mag_io         : inout std_logic ;
    ms_drdy_mag_io        : inout std_logic ;

    magram_clk            : out   std_logic ;
    magram_cs_out         : out   std_logic ;
    magram_mosi_out       : out   std_logic ;
    magram_miso_io        : inout std_logic ;
    magram_writeprot_out  : out   std_logic ;

    mic_clk               : out   std_logic ;
    mic_right_io          : inout std_logic ;
    mic_left_io           : inout std_logic ;

    radio_clk             : out   std_logic ;
    radio_data_io         : inout std_logic_vector (3 downto 0)
  ) ;

end entity Collar ;


architecture structural of Collar is

  --  Establish keep attribute to override optimization removal of signals
  --  needed by SDC files.

  attribute keep              : boolean ;

  --  Master clock information.

  constant master_clk_freq_c  : natural := source_clk_freq_g ;

  signal master_clk           : std_logic ;
  signal master_gated_clk     : std_logic ;
  signal master_gated_inv_clk : std_logic ;
  signal master_gated_en_s    : std_logic ;

  attribute keep of master_gated_en_s   : signal is true ;

  --  Button specifications.

  constant reset_button_c     : natural := 0 ;
  constant sd_start_button_c  : natural := 1 ;

  --  Clock and time signals.

  signal reset_time_bytes     : std_logic_vector (gps_time_bytes_c*8-1
                                                  downto 0) ;
  signal reset_time           : std_logic_vector (gps_time_bits_c-1
                                                  downto 0) ;
  signal gps_time_bytes       : std_logic_vector (gps_time_bytes_c*8-1
                                                  downto 0) ;
  signal gps_time             : std_logic_vector (gps_time_bits_c-1
                                                  downto 0) ;
  signal systime_latch        : std_logic ;
  signal systime_valid        : std_logic ;
  signal systime_vlatch       : std_logic ;
  signal rtc_seconds          : unsigned (epoch70_secbits_c-1 downto 0) ;
  signal rtc_seconds_load     : std_logic ;
  signal rtc_running_seconds  : unsigned (epoch70_secbits_c-1 downto 0) ;
  signal rtc_running_set      : std_logic ;
  signal running_datetime     : std_logic_vector (dt_totalbits_c-1
                                                  downto 0) ;
  signal sunrise_today        : unsigned (epoch70_secbits_c-1 downto 0) ;
  signal sunset_today         : unsigned (epoch70_secbits_c-1 downto 0) ;
  signal sunrise_tomorrow     : unsigned (epoch70_secbits_c-1 downto 0) ;
  signal sunset_tomorrow      : unsigned (epoch70_secbits_c-1 downto 0) ;

  --  Reset information.  The power up signal defaults to zero.

  constant pu_time_c        : real    := 0.5 ;   -- Give sigtap start time.
  constant pu_count_c       : natural :=
              natural (trunc (real (master_clk_freq_c) * pu_time_c)) ;

  signal reset              : std_logic ;
  signal power_up           : std_logic := '0' ;
  signal pu_counter         : unsigned (const_bits (pu_count_c)-1
                                        downto 0) := (others => '0') ;

  constant pb_time_c        : real    := 0.5 ;
  constant pb_count_c       : natural :=
              natural (trunc (real (master_clk_freq_c) * pb_time_c)) ;

  signal reset_pushed       : std_logic := '0' ;
  signal pb_counter         : unsigned (const_bits (pb_count_c)-1
                                        downto 0) := (others => '0') ;

  COMPONENT GlobalClock IS
    PORT
    (
      ena    : IN STD_LOGIC  := '1';
      inclk    : IN STD_LOGIC ;
      outclk    : OUT STD_LOGIC
    );
  END COMPONENT GlobalClock;

  --  Allow JTAG to determine the location code for this executable.

  signal LocationCode       :
            unsigned (const_bits (CP_LocationTbl_c'length-1)-1 downto 0) :=
                TO_UNSIGNED (CP_Loc_code_c,
                             const_bits (CP_LocationTbl_c'length-1)) ;

  attribute noprune                   : boolean ;
  attribute noprune of LocationCode   : signal is true ;

  --  SPI clocks.

  signal spi_clk              : std_logic ;
  signal spi_gated_clk        : std_logic ;
  signal spi_gated_inv_clk    : std_logic ;
  signal spi_gated_en_s       : std_logic ;

  attribute keep of spi_gated_en_s  : signal is true ;

  component GenClock is

    Generic (
      clk_freq_g              : natural   := 10e6 ;
      out_clk_freq_g          : natural   := 1e6 ;
      net_clk_g               : natural   := 0 ;
      net_inv_g               : natural   := 0 ;
      net_gated_g             : natural   := 0 ;
      net_inv_gated_g         : natural   := 0
     ) ;
    Port (
      reset                   : in    std_logic ;
      clk                     : in    std_logic ;
      clk_on_in               : in    std_logic ;
      clk_off_in              : in    std_logic ;
      clk_out                 : out   std_logic ;
      clk_inv_out             : out   std_logic ;
      gated_clk_out           : out   std_logic ;
      gated_clk_inv_out       : out   std_logic
    ) ;

  end component GenClock ;

  --  PC control and status signals.

  signal StatCtlActive          : std_logic ;
  signal PC_StatusSet           : std_logic ;
  signal PC_StatusReg           : std_logic_vector (StatusSignalsCnt_c-1
                                                    downto 0) ;

  alias STAT_BatteryGood        : std_logic is
        PC_StatusReg (StatusSignals'pos (Stat_BatteryGood_e)) ;
  alias STAT_SolarCtlOn       : std_logic is
        PC_StatusReg (StatusSignals'pos (Stat_SolarCtlOn_e)) ;
  alias STAT_SolarCtlMax        : std_logic is
        PC_StatusReg (StatusSignals'pos (Stat_SolarCtlMax_e)) ;
  alias STAT_BattMonLow       : std_logic is
        PC_StatusReg (StatusSignals'pos (Stat_BattMonLow_e)) ;
  alias STAT_ForceStartup       : std_logic is
        PC_StatusReg (StatusSignals'pos (Stat_ForceStartup_e)) ;
  alias STAT_PwrGood2p5       : std_logic is
        PC_StatusReg (StatusSignals'pos (Stat_PwrGood2p5_e)) ;
  alias STAT_PwrGood3p3       : std_logic is
        PC_StatusReg (StatusSignals'pos (Stat_PwrGood3p3_e)) ;


  signal PC_ControlTurnOn       : std_logic_vector (ControlSignalsCnt_c-1
                                                    downto 0) ;

  signal PC_ControlReg          : std_logic_vector (ControlSignalsCnt_c-1
                                                    downto 0) :=
                                      (others => '0') ;

  alias CTL_MainPowerSwitch     : std_logic is
        PC_ControlReg (ControlSignals'pos (Ctl_MainPowerSwitch_e)) ;
  alias CTL_RechargeSwitch      : std_logic is
        PC_ControlReg (ControlSignals'pos (Ctl_RechargeSwitch_e)) ;
  alias CTL_SolarCtlShutdown    : std_logic is
        PC_ControlReg (ControlSignals'pos (Ctl_SolarCtlShutdown_e)) ;
  alias CTL_LevelShifter3p3     : std_logic is
        PC_ControlReg (ControlSignals'pos (Ctl_LevelShifter3p3_e)) ;
  alias CTL_LevelShifter1p8     : std_logic is
        PC_ControlReg (ControlSignals'pos (Ctl_LevelShifter1p8_e)) ;
  alias CTL_InertialOn1p8       : std_logic is
        PC_ControlReg (ControlSignals'pos (Ctl_InertialOn1p8_e)) ;
  alias CTL_InertialOn2p5       : std_logic is
        PC_ControlReg (ControlSignals'pos (Ctl_InertialOn2p5_e)) ;
  alias CTL_MicLeftOn           : std_logic is
        PC_ControlReg (ControlSignals'pos (Ctl_MicLeftOn_e)) ;
  alias CTL_MicRightOn          : std_logic is
        PC_ControlReg (ControlSignals'pos (Ctl_MicRightOn_e)) ;
  alias CTL_SDRAM_On            : std_logic is
        PC_ControlReg (ControlSignals'pos (Ctl_SDRAM_On_e)) ;
  alias CTL_SDCardOn            : std_logic is
        PC_ControlReg (ControlSignals'pos (Ctl_SDCardOn_e)) ;
  alias CTL_MagMemOn            : std_logic is
        PC_ControlReg (ControlSignals'pos (Ctl_MagMemOn_e)) ;
  alias CTL_GPS_On              : std_logic is
        PC_ControlReg (ControlSignals'pos (Ctl_GPS_On_e)) ;
  alias CTL_DataTX_On           : std_logic is
        PC_ControlReg (ControlSignals'pos (Ctl_DataTX_On_e)) ;
  alias CTL_FPGA_Shutdown       : std_logic is
        PC_ControlReg (ControlSignals'pos (Ctl_FPGA_Shutdown_e)) ;
  alias CTL_FLASH_Granted       : std_logic is
        PC_ControlReg (ControlSignals'pos (Ctl_FLASH_Granted_e)) ;

  --  Memory resouce sharing constants and signals.
  --  Memory sharing involves each component sharing a memory bus, building
  --  a vector that is a concatination of all its control and output data
  --  signals.  This vector is added to a table of vectors for all
  --  components that share the memory bus.  Resource allocation is used
  --  to determine the current bus user and its control vector is mapped
  --  to the memory bus.
  --  When a component does not write to memory it uses the 'none'
  --  constants for that part of the combined signal.

  --  Shared GPS Memory constants and signals.

  constant gpsmem_bytecnt_c     : natural := 1024 ;
  constant gpsmem_databits_c    : natural := 8 ;
  constant gpsmem_elementcnt_c  : natural := 8 * gpsmem_bytecnt_c /
                                                 gpsmem_databits_c ;

  constant gpsmem_addrbits_c    : natural :=
                                      const_bits (gpsmem_elementcnt_c-1) ;
  constant gpsmem_rdwr_enbits_c : natural := 2 ;
  constant gpsmem_clkbits_c     : natural := 1 ;
  constant gpsmem_iobits_c      : natural := gpsmem_databits_c +
                                             gpsmem_addrbits_c +
                                             gpsmem_rdwr_enbits_c +
                                             gpsmem_clkbits_c ;

  constant gpsmem_wrto_none_c   : std_logic_vector (gpsmem_databits_c-1
                                                    downto 0) :=
                                                        (others => '0') ;
  constant gpsmem_wren_none_c   : std_logic := '0' ;

  --  Memory requestors.

  constant gpsmemrq_flashblk_c    : natural := 0 ;
  constant gpsmemrq_systemtime_c  : natural := gpsmemrq_flashblk_c    + 1 ;

  constant gpsmemrq_count_c       : natural := gpsmemrq_systemtime_c  + 1 ;

  signal gpsmem_requesters        : std_logic_vector (gpsmemrq_count_c-1
                                                      downto 0) ;
  signal gpsmem_receivers         : std_logic_vector (gpsmemrq_count_c-1
                                                      downto 0) ;

  signal gpsmem_input_tbl         : std_logic_2D (gpsmemrq_count_c-1
                                                  downto 0,
                                                  gpsmem_iobits_c-1
                                                  downto 0) ;

  signal gpsmemdst_readfrom       : std_logic_vector (gpsmem_databits_c-1
                                                      downto 0) ;

  --------------------------------------------------------------------------
  --  Shared Magnetic Memory constants and signals.
  --------------------------------------------------------------------------

  constant magmem_bytecnt_c     : natural := magmem_buffer_bytes ;
  constant magmem_databits_c    : natural := 8 * magmem_data_width_a_bytes ;
  constant magmem_elementcnt_c  : natural := 8 * magmem_bytecnt_c /
                                                 magmem_databits_c ;

  constant magmem_addrbits_c    : natural :=
                                      const_bits (magmem_elementcnt_c-1) ;
  constant magmem_rdwr_enbits_c : natural := 2 ;
  constant magmem_clkbits_c     : natural := 1 ;
  constant magmem_iobits_c      : natural := magmem_databits_c +
                                             magmem_addrbits_c +
                                             magmem_rdwr_enbits_c +
                                             magmem_clkbits_c  ;

  constant magmem_wrto_none_c   : std_logic_vector (magmem_databits_c-1
                                                    downto 0) :=
                                                        (others => '0') ;
  constant magmem_wren_none_c   : std_logic := '0' ;

  --  Memory requestors.

  constant magmemrq_magmem_c    : natural := 0 ;
  constant magmemrq_flashblk_c  : natural := magmemrq_magmem_c      + 1 ;
  constant magmemrq_sdcard_c    : natural := magmemrq_flashblk_c    + 1 ;

  constant magmemrq_count_c     : natural := magmemrq_sdcard_c      + 1 ;

  signal magmem_requesters      : std_logic_vector (magmemrq_count_c-1
                                                    downto 0) ;
  signal magmem_receivers       : std_logic_vector (magmemrq_count_c-1
                                                    downto 0) ;

  signal magmem_input_tbl       : std_logic_2D (magmemrq_count_c-1 downto 0,
                                                magmem_iobits_c-1 downto 0) ;

  signal magmemsrc_readfrom     : std_logic_vector (magmem_databits_c-1
                                                    downto 0) ;

  --------------------------------------------------------------------------
  --  Event Logging memory constants and signals.
  --------------------------------------------------------------------------

  constant eventcnt_events_c    : natural := collar_event_cnt_c ;

  constant eventcnt_countbits_c : natural := 8 ;

  constant eventcnt_membytes_c  : natural := 1024 ;

  constant eventcnt_bytes_c     : natural :=
              natural (trunc (real ((eventcnt_events_c - 1)*
                                    eventcnt_countbits_c) / 8.0)) + 1 ;

  constant eventcnt_databits_c  : natural := eventcnt_countbits_c ;
  constant eventcnt_addrbits_c  : natural :=
              const_bits (eventcnt_membytes_c * 8 /
                          eventcnt_databits_c - 1) ;

  signal evmemdst_clk           : std_logic ;
  signal evmemdst_readfrom      : std_logic_vector (eventcnt_databits_c-1
                                                    downto 0) ;
  signal evmemdst_writeto       : std_logic_vector (eventcnt_databits_c-1
                                                    downto 0) ;
  signal evmemdst_addr          : std_logic_vector (eventcnt_addrbits_c-1
                                                    downto 0) ;
  signal evmemdst_read_en       : std_logic ;
  signal evmemdst_write_en      : std_logic ;

  --  Event increment vector signals.

  signal eventcnt_clear         : std_logic ;
  signal eventcnt_lock          : std_logic ;
  signal eventcnt_changed       : std_logic ;
  signal eventcnt_busy          : std_logic ;

  signal eventcnt_incr          : std_logic_vector (eventcnt_events_c-1
                                                    downto 0) ;

  alias ev_MainPowerSwitchOn    : std_logic is
          eventcnt_incr (Collar_Events'pos (CE_MainPowerSwitchOn_e)) ;
  alias ev_MainPowerSwitchOff   : std_logic is
          eventcnt_incr (Collar_Events'pos (CE_MainPowerSwitchOff_e)) ;
  alias ev_RechargeSwitchOn   : std_logic is
          eventcnt_incr (Collar_Events'pos (CE_RechargeSwitchOn_e)) ;
  alias ev_RechargeSwitchOff    : std_logic is
          eventcnt_incr (Collar_Events'pos (CE_RechargeSwitchOff_e)) ;
  alias ev_SolarCtlShutdownOn   : std_logic is
          eventcnt_incr (Collar_Events'pos (CE_SolarCtlShutdownOn_e)) ;
  alias ev_SolarCtlShutdownOff    : std_logic is
          eventcnt_incr (Collar_Events'pos (CE_SolarCtlShutdownOff_e)) ;
  alias ev_LevelShifter3p3On    : std_logic is
          eventcnt_incr (Collar_Events'pos (CE_LevelShifter3p3On_e)) ;
  alias ev_LevelShifter3p3Off   : std_logic is
          eventcnt_incr (Collar_Events'pos (CE_LevelShifter3p3Off_e)) ;
  alias ev_LevelShifter1p8On    : std_logic is
          eventcnt_incr (Collar_Events'pos (CE_LevelShifter1p8On_e)) ;
  alias ev_LevelShifter1p8Off   : std_logic is
          eventcnt_incr (Collar_Events'pos (CE_LevelShifter1p8Off_e)) ;
  alias ev_InertialOn1p8    : std_logic is
          eventcnt_incr (Collar_Events'pos (CE_InertialOn1p8_e)) ;
  alias ev_InertialOff2p5   : std_logic is
          eventcnt_incr (Collar_Events'pos (CE_InertialOff2p5_e)) ;
  alias ev_MicLeftOn    : std_logic is
          eventcnt_incr (Collar_Events'pos (CE_MicLeftOn_e)) ;
  alias ev_MicLeftOff   : std_logic is
          eventcnt_incr (Collar_Events'pos (CE_MicLeftOff_e)) ;
  alias ev_MicRightOn   : std_logic is
          eventcnt_incr (Collar_Events'pos (CE_MicRightOn_e)) ;
  alias ev_MicRightOff    : std_logic is
          eventcnt_incr (Collar_Events'pos (CE_MicRightOff_e)) ;
  alias ev_SDRAM_On   : std_logic is
          eventcnt_incr (Collar_Events'pos (CE_SDRAM_On_e)) ;
  alias ev_SDRAM_Off    : std_logic is
          eventcnt_incr (Collar_Events'pos (CE_SDRAM_Off_e)) ;
  alias ev_SDCardOn   : std_logic is
          eventcnt_incr (Collar_Events'pos (CE_SDCardOn_e)) ;
  alias ev_SDCardOff    : std_logic is
          eventcnt_incr (Collar_Events'pos (CE_SDCardOff_e)) ;
  alias ev_GPS_On   : std_logic is
          eventcnt_incr (Collar_Events'pos (CE_GPS_On_e)) ;
  alias ev_GPS_Off    : std_logic is
          eventcnt_incr (Collar_Events'pos (CE_GPS_Off_e)) ;
  alias ev_DataTX_On    : std_logic is
          eventcnt_incr (Collar_Events'pos (CE_DataTX_On_e)) ;
  alias ev_DataTX_Off   : std_logic is
          eventcnt_incr (Collar_Events'pos (CE_DataTX_Off_e)) ;
  alias ev_BatteryGoodOn    : std_logic is
          eventcnt_incr (Collar_Events'pos (CE_BatteryGoodOn_e)) ;
  alias ev_BatteryGoodOff   : std_logic is
          eventcnt_incr (Collar_Events'pos (CE_BatteryGoodOff_e)) ;
  alias ev_SolarCtlOn   : std_logic is
          eventcnt_incr (Collar_Events'pos (CE_SolarCtlOn_e)) ;
  alias ev_SolarCtlOff    : std_logic is
          eventcnt_incr (Collar_Events'pos (CE_SolarCtlOff_e)) ;
  alias ev_BattMonLowOn   : std_logic is
          eventcnt_incr (Collar_Events'pos (CE_BattMonLowOn_e)) ;
  alias ev_BattMonLowOff    : std_logic is
          eventcnt_incr (Collar_Events'pos (CE_BattMonLowOff_e)) ;
  alias ev_ForceStartupOn   : std_logic is
          eventcnt_incr (Collar_Events'pos (CE_ForceStartupOn_e)) ;
  alias ev_ForceStartupOff    : std_logic is
          eventcnt_incr (Collar_Events'pos (CE_ForceStartupOff_e)) ;
  alias ev_PwrGood2p5On   : std_logic is
          eventcnt_incr (Collar_Events'pos (CE_PwrGood2p5On_e)) ;
  alias ev_PwrGood2p5Off    : std_logic is
          eventcnt_incr (Collar_Events'pos (CE_PwrGood2p5Off_e)) ;
  alias ev_PwrGood3p3On   : std_logic is
          eventcnt_incr (Collar_Events'pos (CE_PwrGood3p3On_e)) ;
  alias ev_PwrGood3p3Off    : std_logic is
          eventcnt_incr (Collar_Events'pos (CE_PwrGood3p3Off_e)) ;

  --------------------------------------------------------------------------
  --  SDRAM constants and signals.
  --------------------------------------------------------------------------

  constant sdram_rowbytes_c     : natural := sdram_space_g.ROWBITS / 8 ;

  constant sdram_bytes_c        : natural := sdram_space_g.BANKS *
                                             sdram_space_g.ROWCOUNT *
                                             sdram_rowbytes_c ;

  constant outmem_bytecnt_c     : natural := 4096 ;
  constant outmem_rdwidth_c     : natural := 8 ;

  constant outmem_buffrows_c    : natural := 1 ;
  constant outmem_buffcount_c   : natural :=
              outmem_bytecnt_c / (sdram_rowbytes_c * outmem_buffrows_c) ;

  constant outmem_rdelements_c  : natural :=
              8 * outmem_bytecnt_c / outmem_rdwidth_c ;

  constant outmem_rdaddrbits_c  : natural :=
              const_bits (outmem_rdelements_c - 1) ;

  constant inmem_bytecnt_c      : natural := 4096 ;
  constant inmem_wrwidth_c      : natural := 8 ;

  constant inmem_buffouts_c     : natural := 1 ;
  constant inmem_buffcount_c    : natural :=
              inmem_bytecnt_c / (sdram_rowbytes_c * outmem_buffrows_c *
                                 inmem_buffouts_c) ;

  constant inmem_wrelements_c   : natural :=
              8 * inmem_bytecnt_c / inmem_wrwidth_c ;

  constant inmem_wraddrbits_c   : natural :=
              const_bits (inmem_wrelements_c - 1) ;

  signal sdram_ready            : std_logic ;
  signal sdram_empty            : std_logic ;
  signal sdram_forceout         : std_logic ;

  signal sdram_inready          : std_logic ;
  signal sdram_inwr_data        : std_logic_vector (inmem_wrwidth_c-1
                                                    downto 0) ;
  signal sdram_inwr_addr        : std_logic_vector (inmem_wraddrbits_c-1
                                                    downto 0) ;
  signal sdram_inwr_en          : std_logic ;
  signal sdram_inwr_clk         : std_logic ;

  signal sdram_outready         : std_logic ;
  signal sdram_outwriting       : std_logic ;
  signal sdram_outamt           : unsigned (const_bits (sdram_bytes_c-1)-1
                                            downto 0) ;
  signal sdram_outrd_data       : std_logic_vector (outmem_rdwidth_c-1
                                                    downto 0) ;
  signal sdram_outrd_addr       : std_logic_vector (outmem_rdaddrbits_c-1
                                                    downto 0) ;
  signal sdram_outrd_en         : std_logic ;
  signal sdram_outrd_clk        : std_logic ;

  --------------------------------------------------------------------------
  --  SD Card constants and signals.
  --------------------------------------------------------------------------

  constant sdcard_blksize_c     : natural := 512 ;
  constant sdcard_blknobits_c   : natural := 32 ;

  signal sdcard_start           : std_logic ;

  signal sdcard_critdone        : std_logic ;
  signal sdcard_critpast        : std_logic_vector (7 downto 0) ;

  --------------------------------------------------------------------------
  --  GPS signals.
  --------------------------------------------------------------------------

  signal gps_init               : std_logic ;
  signal gps_ready              : std_logic ;

  signal gps_databanks          : std_logic_vector (msg_ram_blocks_c-1
                                                    downto 0) ;
  signal aop_running            : std_logic ;

  --  GPS dual port RAM communication signals.

  constant gpsmemsrc_addrbits_c : natural := gpsmem_addrbits_c ;
  constant gpsmemsrc_databits_c : natural := gpsmem_databits_c ;

  signal gpsmemsrc_addr         : std_logic_vector (gpsmemsrc_addrbits_c-1
                                                    downto 0) ;
  signal gpsmemsrc_clk          : std_logic ;
  signal gpsmemsrc_writeto      : std_logic_vector (gpsmemsrc_databits_c-1
                                                    downto 0) ;
  signal gpsmemsrc_readfrom     : std_logic_vector (gpsmemsrc_databits_c-1
                                                    downto 0) ;
  signal gpsmemsrc_read_en      : std_logic ;
  signal gpsmemsrc_write_en     : std_logic ;

  --------------------------------------------------------------------------
  --  Magnetic Memory dual port RAM communication signals.
  --------------------------------------------------------------------------

  signal magmemdst_addr         : std_logic_vector (magmem_addrbits_c-1
                                                    downto 0) ;
  signal magmemdst_readfrom     : std_logic_vector (magmem_databits_c-1
                                                    downto 0) ;
  signal magmemdst_writeto      : std_logic_vector (magmem_databits_c-1
                                                    downto 0) ;
  signal magmemdst_read_en      : std_logic ;
  signal magmemdst_write_en     : std_logic ;
  signal magmemdst_clk          : std_logic ;

  signal magmem_buff_busy       : std_logic ;

  --------------------------------------------------------------------------
  --  Inertial module constants and signals.
  --------------------------------------------------------------------------

  constant im_datalen_c     : natural := 2 ;
  constant im_databits_c    : natural := im_datalen_c * 8 ;

  signal im_startup         : std_logic ;
  signal im_startup_done    : std_logic ;
  signal im_gyro_data_rdy   : std_logic ;
  signal im_accel_data_rdy  : std_logic ;
  signal im_mag_data_rdy    : std_logic ;
  signal im_temp_data_rdy   : std_logic ;
  signal im_gyro_data_x     : std_logic_vector (im_databits_c-1 downto 0) ;
  signal im_gyro_data_y     : std_logic_vector (im_databits_c-1 downto 0) ;
  signal im_gyro_data_z     : std_logic_vector (im_databits_c-1 downto 0) ;
  signal im_accel_data_x    : std_logic_vector (im_databits_c-1 downto 0) ;
  signal im_accel_data_y    : std_logic_vector (im_databits_c-1 downto 0) ;
  signal im_accel_data_z    : std_logic_vector (im_databits_c-1 downto 0) ;
  signal im_mag_data_x      : std_logic_vector (im_databits_c-1 downto 0) ;
  signal im_mag_data_y      : std_logic_vector (im_databits_c-1 downto 0) ;
  signal im_mag_data_z      : std_logic_vector (im_databits_c-1 downto 0) ;
  signal im_temp_data       : std_logic_vector (im_databits_c-1 downto 0) ;
  signal im_gyro_time       : std_logic_vector (gps_time_bytes_c*8-1
                                                downto 0) ;
  signal im_accel_time      : std_logic_vector (gps_time_bytes_c*8-1
                                                downto 0) ;
  signal im_mag_time        : std_logic_vector (gps_time_bytes_c*8-1
                                                downto 0) ;
  signal im_temp_time       : std_logic_vector (gps_time_bytes_c*8-1
                                                downto 0) ;

  --------------------------------------------------------------------------
  --  Magnetic memory constants and signals.
  --------------------------------------------------------------------------

  constant mm_buffbytes_c   : natural := magmem_bytecnt_c ;
  constant mm_buffnum_c     : natural := magmem_buffer_num ;

  signal mm_startup         : std_logic ;
  signal mm_startup_done    : std_logic ;
  signal mm_buffno          : std_logic_vector (
                                    const_bits (mm_buffnum_c-1)-1 downto 0) ;

  --------------------------------------------------------------------------
  --  Microphone constants and signals.
  --------------------------------------------------------------------------

  constant mic_sample_bits_c  : natural := 16 ;
  constant mic_sample_bytes_c : natural :=
              natural (trunc (real (mic_sample_bits_c - 1) / 8.0)) + 1 ;

  signal mic_right_sample     : std_logic_vector (mic_sample_bits_c-1
                                                  downto 0) ;
  signal mic_right_sample_clk : std_logic ;

  signal mic_left_sample      : std_logic_vector (mic_sample_bits_c-1
                                                  downto 0) ;
  signal mic_left_sample_clk  : std_logic ;

  --------------------------------------------------------------------------
  --  Real-time Clock constants and signals.
  --------------------------------------------------------------------------

  --constant rtc_time_bytes_c   : natural := epoch70_secbits_c / 8 ;

  constant rtc_time_bytes_c   : natural := 4 ;
  
  constant tod_bytes : natural := 4;
  constant alarm_bytes : natural := 3;

  signal rtc_time             : std_logic_vector (rtc_time_bytes_c*8-1
                                                  downto 0) :=
                                                      (others => '0') ;
                                                      
                                                      
             
  signal    tod_set_signal          :     std_logic := '0';
  signal    tod_set_done_signal     :     std_logic := '0';
  signal    tod_set             :     std_logic_vector(tod_bytes*8-1 downto 0);
    
    
  signal    tod_get_signal        :    std_logic := '0';
  signal    tod_signal            :    std_logic_vector(tod_bytes*8-1 downto 0);     
  signal    tod_get_valid_signal  :    std_logic := '0';

  signal    alarm_set_signal          :     std_logic := '0';    
  signal    alarm_signal              :     std_logic_vector(alarm_bytes*8-1 downto 0);
  signal    alarm_set_done_signal     :     std_logic := '0';
  
  
  signal    rtc_interrupt_enable_signal :   std_logic;
  
  
  signal rtc_startup        : std_logic;  
  signal rtc_startup_done   : std_logic;
  
  
  --------------------------------------------------------------------------
  --  Battery Monitor Inupts/Ouputs
  --------------------------------------------------------------------------
  
  
  signal batmon_startup: std_logic;
  
  signal rem_cap_mah_signal : std_logic_vector (15 downto 0);
  signal inst_cur_ma_signal : std_logic_vector (15 downto 0);
  signal voltage_mv_signal : std_logic_vector (15 downto 0);
  
  signal voltage_mv_valid_signal : std_logic;
  signal inst_cur_ma_valid_signal : std_logic;
  signal rem_cap_mah_valid_signal : std_logic;


  --------------------------------------------------------------------------
  --  Constants and signals to control logging of information to the SDCard.
  --  The logging sequence number is started beyond its last known value
  --  when logging begins after a restart.
  --  Status information can be logged by force.
  --  All buffered data can be flushed to the SDCard.
  --------------------------------------------------------------------------

  constant SDLogging_seqbits_c  : natural := 32 ;

  signal SDLogging_seqno        : std_logic_vector (SDLogging_seqbits_c-1
                                                    downto 0) :=
                                                        (others => '0') ;

  signal SDLogging_status       : std_logic := '0' ;
  signal SDLogging_flush        : std_logic := '0' ;

  component Startup_Shutdown is
    Generic (
      clk_freq_g            : natural := 50e6
    );
    Port (
      clk                 : in    std_logic ;
      rst_n               : in    std_logic ;
      pc_control_reg_out  : out std_logic_vector (ControlSignalsCnt_c-1
                                            downto 0);     
      pc_control_reg_in  : in   std_logic_vector (ControlSignalsCnt_c-1
                                                  downto 0) ;                                           
      pc_status_set_in          : in      std_logic;
      sd_contr_start_out        : out   std_logic ;       
      sd_contr_done_in          : in    std_logic ;   
      sdram_start_out           : out   std_logic ;
      sdram_done_in             : in    std_logic ;
      imu_start_out             : out   std_logic ;
      imu_done_in               : in    std_logic ;
      rtc_start_out             : out   std_logic ;
      rtc_done_in               : in    std_logic ;
      batmon_start_out          : out   std_logic ;
      batmon_done_in            : in    std_logic ;
      mems_start_out            : out   std_logic ;
      mems_done_in              : in    std_logic ;
      mag_start_out             : out   std_logic ;
      mag_done_in               : in    std_logic ;
      gps_start_out             : out   std_logic ;
      gps_done_in               : in    std_logic ;
      txrx_start_out            : out   std_logic ;
      txrx_done_in              : in    std_logic ;
      shutdown_in               : in    std_logic ;
      statctl_startup_out       : out   std_logic;
      rem_cap_mah_valid_in      : in    std_logic ; 
      rem_cap_mah_in            : in    std_logic_vector (15 downto 0)
  ) ;
  
    end component Startup_Shutdown ;

begin

  --------------------------------------------------------------------------
  --  Startup Machine
  --  System startup sequencing and setting of the control register.
  --------------------------------------------------------------------------

  
  signal shutdown_master           :  std_logic := '0';
  signal statctl_startup_signal    :  std_logic;
  
  
  i_startup_0 : Startup_Shutdown
    Generic Map (
      clk_freq_g              => spi_clk_freq_c
    )
    Port Map(
      clk                 => spi_clk,
      rst_n               => not reset,
      
      pc_control_reg_out        =>  PC_ControlReg,   
      pc_control_reg_in         =>  PC_ControlReg_signal,        
      pc_status_set_in          =>  PC_StatusSet,
      sd_contr_start_out        =>  sdcard_start,
      sd_contr_done_in          =>  '1',
      --sdram_start_out             : out  std_logic ;
      sdram_done_in             => sdram_ready,
      imu_start_out             => im_startup,
      imu_done_in               => im_startup_done,
      rtc_start_out             => rtc_startup,
      rtc_done_in               => rtc_startup_done,
      batmon_start_out          => batmon_startup,
      batmon_done_in            => '1',
      --mems_start_out            : out std_logic ;
      mems_done_in              => '1',
      mag_start_out             => mm_startup,
      mag_done_in               => mm_startup_done,
      --gps_start_out             : out   std_logic ;
      gps_done_in               => '1',
      --txrx_start_out            : out   std_logic ;
      txrx_done_in              => '1',
      shutdown_in               => shutdown_master,
      statctl_startup_out       => statctl_startup_signal,
      rem_cap_mah_valid_in      => rem_cap_mah_valid_signal,
      rem_cap_mah_in            => rem_cap_mah_signal
      

    ) ;

  PC_ControlReg                 <= PC_ControlReg or PC_ControlTurnOn ;


  --------------------------------------------------------------------------
  --  SPI clock.
  --  The gated clock is turned on when a component that needs it becomes
  --  active.
  --  NOTE: Gate turn-on takes over one source clock cycles to complete.
  --        As this is shorter than one half SPI clock cycle it is not a
  --        problem.  If a faster response time is needed then another
  --        mechanism must be used.
  --------------------------------------------------------------------------

  spi_clock : GenClock
    Generic Map (
      clk_freq_g              => master_clk_freq_c,
      out_clk_freq_g          => spi_clk_freq_c,
      net_clk_g               => 1,
      net_gated_g             => 1,
      net_inv_gated_g         => 0
    )
    Port Map (
      reset                   => reset,
      clk                     => master_clk,
      clk_on_in               => spi_gated_en_s,
      clk_off_in              => not spi_gated_en_s,
      clk_out                 => spi_clk,
      gated_clk_out           => spi_gated_clk,
      gated_clk_inv_out       => spi_gated_inv_clk
    ) ;

  spi_gated_en_s        <= StatCtlActive                           or
                           magmem_requesters (magmemrq_magmem_c)   or
                           magmem_receivers  (magmemrq_magmem_c)   or
                           magmem_requesters (magmemrq_flashblk_c) or
                           magmem_receivers  (magmemrq_flashblk_c) or
                           gpsmem_requesters (gpsmemrq_flashblk_c) or
                           gpsmem_receivers  (gpsmemrq_flashblk_c) ;


  --------------------------------------------------------------------------
  --  Master clock.
  --  The gated clock is turned on when the shared gps memory port is used
  --  and under other conditions.
  --------------------------------------------------------------------------

  master_clock : GenClock
    Generic Map (
      clk_freq_g              => master_clk_freq_c,
      out_clk_freq_g          => master_clk_freq_c,
      net_clk_g               => 1,
      net_gated_g             => 1,
      net_inv_gated_g         => 1
    )
    Port Map (
      reset                   => '0',
      clk                     => source_clk,
      clk_on_in               => master_gated_en_s,
      clk_off_in              => not master_gated_en_s,
      clk_out                 => master_clk,
      gated_clk_out           => master_gated_clk,
      gated_clk_inv_out       => master_gated_inv_clk
    ) ;

  master_gated_en_s     <= '1' when ((unsigned (gpsmem_requesters) /= 0)  or
                                     (unsigned (gpsmem_receivers)  /= 0)  or
                                     eventcnt_busy    = '1'               or
                                     magmem_buff_busy = '1')
                               else '0' ;


  --------------------------------------------------------------------------
  --  System Time clocks.
  --------------------------------------------------------------------------

  use_StrClk:
    if (Collar_Control_useStrClk_c = '1') generate

      component SystemTime is
        Generic (
          clk_freq_g          : natural := 50e3 ;
          gpsmem_addrbits_g   : natural := 10 ;
          gpsmem_databits_g   : natural :=  8 ;
          timezone_g          : integer := -7 * 60 * 60 ;
          dst_start_mth_g     : natural :=  3 ;
          dst_start_day_g     : natural :=  8 ;
          dst_start_hr_g      : natural :=  2 ;
          dst_start_min_g     : natural :=  0 ;
          dst_end_mth_g       : natural := 11 ;
          dst_end_day_g       : natural :=  1 ;
          dst_end_hr_g        : natural :=  2 ;
          dst_end_min_g       : natural :=  0 ;
          dst_seconds_g       : natural := 60 * 60
        ) ;
        Port (
          reset               : in    std_logic ;
          clk                 : in    std_logic ;
          startup_time_out    : out   std_logic_vector (gps_time_bits_c-1
                                                        downto 0) ;
          startup_bytes_out   : out   std_logic_vector (gps_time_bytes_c*8-1
                                                        downto 0) ;
          gps_time_out        : out   std_logic_vector (gps_time_bits_c-1
                                                        downto 0) ;
          gps_bytes_out       : out   std_logic_vector (gps_time_bytes_c*8-1
                                                        downto 0) ;

          rtc_sec_in          : in    unsigned (epoch70_secbits_c-1 downto 0) ;
          rtc_sec_load_in     : in    std_logic ;
          rtc_sec_out         : out   unsigned (epoch70_secbits_c-1 downto 0) ;
          rtc_sec_set_out     : out   std_logic ;
          rtc_datetime_out    : out   std_logic_vector (dt_totalbits_c-1
                                                        downto 0) ;

          time_latch_out      : out   std_logic ;
          time_valid_out      : out   std_logic ;
          valid_latch_out     : out   std_logic ;

          gpsmem_tmbank_in    : in    std_logic ;
          gpsmem_req_out      : out   std_logic ;
          gpsmem_rcv_in       : in    std_logic ;
          gpsmem_addr_out     : out   std_logic_vector (gpsmem_addrbits_g-1
                                                        downto 0) ;
          gpsmem_datafrom_in  : in    std_logic_vector (gpsmem_databits_g-1
                                                        downto 0) ;
          gpsmem_readen_out   : out   std_logic ;

          alarm_time_in       : in    std_logic_vector (dt_totalbits_c-1
                                                        downto 0) ;
          alarm_time_out      : out   unsigned  (epoch70_secbits_c-1 downto 0)
        ) ;
      end component SystemTime ;

      --  System Time to GPS Memory communications signals.

      signal st_gpsmem_clk      : std_logic ;
      signal st_gpsmem_rd_en    : std_logic ;
      signal st_gpsmem_addr     : std_logic_vector (gpsmem_addrbits_c-1
                                                    downto 0) ;
      signal st_gpsmem_control  : std_logic_vector (gpsmem_iobits_c-1
                                                      downto 0) ;

      --  Sunrise/Sunset signals.

      signal noon_datetime        : std_logic_vector (dt_totalbits_c-1
                                                      downto 0) ;
      signal noon_seconds         : unsigned (epoch70_secbits_c-1 downto 0) ;

      signal sunrise_today_out    : unsigned (epoch70_secbits_c-1 downto 0) ;
      signal sunset_today_out     : unsigned (epoch70_secbits_c-1 downto 0) ;
      signal sunrise_tomorrow_out : unsigned (epoch70_secbits_c-1 downto 0) ;
      signal sunset_tomorrow_out  : unsigned (epoch70_secbits_c-1 downto 0) ;

      component SunriseSunset is
        Generic (
          location_code_g       : natural :=  0 ;
          longitude_g           : real    := -111.0525791 ;
          timezone_g            : integer := -7 * 60 * 60 ;
          dst_offset_g          : integer := 60 * 60
        ) ;
        Port (
          reset                 : in    std_logic ;
          rtc_sec_in            : in    unsigned (epoch70_secbits_c-1 downto 0) ;
          rtc_datetime_in       : in    std_logic_vector (dt_totalbits_c-1
                                                          downto 0) ;
          alarm_time_out        : out   std_logic_vector (dt_totalbits_c-1
                                                          downto 0) ;
          alarm_time_in         : in    unsigned (epoch70_secbits_c-1 downto 0) ;
          sunrise_today_out     : out   unsigned (epoch70_secbits_c-1 downto 0) ;
          sunset_today_out      : out   unsigned (epoch70_secbits_c-1 downto 0) ;
          sunrise_tomorrow_out  : out   unsigned (epoch70_secbits_c-1 downto 0) ;
          sunset_tomorrow_out   : out   unsigned (epoch70_secbits_c-1 downto 0)
        ) ;
      end component SunriseSunset ;

    begin

      system_clock : SystemTime
        Generic Map (
          clk_freq_g          => master_clk_freq_c,
          gpsmem_addrbits_g   => gpsmem_addrbits_c,
          gpsmem_databits_g   => gpsmem_databits_c,
          timezone_g          => CP_CurrentLocation_c.timezone,
          dst_start_mth_g     => CP_CurrentLocation_c.dst_start_month,
          dst_start_day_g     => CP_CurrentLocation_c.dst_start_mday,
          dst_start_hr_g      => CP_CurrentLocation_c.dst_start_hour,
          dst_start_min_g     => CP_CurrentLocation_c.dst_start_minute,
          dst_end_mth_g       => CP_CurrentLocation_c.dst_end_month,
          dst_end_day_g       => CP_CurrentLocation_c.dst_end_mday,
          dst_end_hr_g        => CP_CurrentLocation_c.dst_end_hour,
          dst_end_min_g       => CP_CurrentLocation_c.dst_end_minute,
          dst_seconds_g       => CP_CurrentLocation_c.dst_change
        )
        Port Map (
          reset               => reset,
          clk                 => master_clk,
          startup_time_out    => reset_time,
          startup_bytes_out   => reset_time_bytes,
          gps_time_out        => gps_time,
          gps_bytes_out       => gps_time_bytes,
          rtc_sec_in          => rtc_seconds,
          rtc_sec_load_in     => rtc_seconds_load,
          rtc_sec_out         => rtc_running_seconds,
          rtc_sec_set_out     => rtc_running_set,
          rtc_datetime_out    => running_datetime,
          time_latch_out      => systime_latch,
          time_valid_out      => systime_valid,
          valid_latch_out     => systime_vlatch,
          gpsmem_tmbank_in    => gps_databanks (msg_ubx_tim_tm2_ramblock_c),
          gpsmem_req_out      => gpsmem_requesters (gpsmemrq_systemtime_c),
          gpsmem_rcv_in       => gpsmem_receivers  (gpsmemrq_systemtime_c),
          gpsmem_addr_out     => st_gpsmem_addr,
          gpsmem_datafrom_in  => gpsmemdst_readfrom,
          gpsmem_readen_out   => st_gpsmem_rd_en,
          alarm_time_in       => noon_datetime,
          alarm_time_out      => noon_seconds
        ) ;

      st_gpsmem_clk       <= master_gated_inv_clk ;

      st_gpsmem_control   <= st_gpsmem_clk        &
                             gpsmem_wren_none_c   & st_gpsmem_rd_en   &
                             gpsmem_wrto_none_c   & st_gpsmem_addr ;

      set2D_element (gpsmemrq_systemtime_c, st_gpsmem_control,
                     gpsmem_input_tbl) ;

      --  Calculate the sunrise/sunset times.

      sunrise_set : SunriseSunset
        Generic Map (
          location_code_g       => CP_Loc_Code_c,
          longitude_g           => CP_CurrentLocation_c.longitude,
          timezone_g            => CP_CurrentLocation_c.timezone,
          dst_offset_g          => CP_CurrentLocation_c.dst_change
        )
        Port Map (
          reset                 => reset,
          rtc_sec_in            => rtc_running_seconds,
          rtc_datetime_in       => running_datetime,
          alarm_time_out        => noon_datetime,
          alarm_time_in         => noon_seconds,
          sunrise_today_out     => sunrise_today,
          sunset_today_out      => sunset_today,
          sunrise_tomorrow_out  => sunrise_tomorrow,
          sunset_tomorrow_out   => sunset_tomorrow
        ) ;

  end generate use_StrClk ;

  --------------------------------------------------------------------------
  --  I2C bus.
  --------------------------------------------------------------------------

  no_use_I2C:
    if (Collar_Control_useI2C_c = '0') generate

      i2c_clk_io              <= 'Z' ;
      i2c_data_io             <= 'Z' ;

    end generate no_use_I2C ;

  --------------------------------------------------------------------------
  --  Power Controller.
  --------------------------------------------------------------------------

  --  Power Controller SPI communications channel.

  use_PC:
    if (Collar_Control_usePC_c = '1') generate

      component StatCtlSPI_FPGA is
        Generic (
          status_bits_g           : natural := 16 ;
          control_bits_g          : natural := 16 ;
          flash_bytes_transfer    : natural := 0 ;
          data_length_bit_width_g : natural := 8
        ) ;
        Port (
          clk                     : in    std_logic ;
          rst_n                   : in    std_logic ;
          status_out              : out   std_logic_vector (status_bits_g-1
                                                            downto 0) ;
          status_chg_in           : in    std_logic ;
          status_set_out          : out   std_logic ;
          control_in              : in    std_logic_vector (control_bits_g-1
                                                            downto 0) ;
          busy_out                : out   std_logic ;
          
          startup_in              : in    std_logic;

          sclk                    : out   std_logic ;
          mosi                    : out   std_logic ;
          miso                    : in    std_logic ;
          cs_n                    : out   std_logic
        ) ;
      end component StatCtlSPI_FPGA ;

      --  Signals for activating communications.

      signal PC_ControlRegLast    : std_logic_vector (PC_ControlReg'length-1
                                                      downto 0) :=
                                                          (others => '0') ;

    begin

      pc_spi : StatCtlSPI_FPGA
        Generic Map (
          status_bits_g               => StatusSignalsCnt_c,
          control_bits_g              => ControlSignalsCnt_c,
          flash_bytes_transfer        => 0,
          data_length_bit_width_g     => 8
        )
        Port Map (
          clk                         => spi_gated_clk,
          rst_n                       => not reset,
          status_out                  => PC_StatusReg,
          status_chg_in               => pc_statchg_in,
          status_set_out              => PC_StatusSet,
          control_in                  => PC_ControlReg,
          busy_out                    => StatCtlActive,
          startup_in                  => statctl_startup_signal,

          sclk                        => pc_spi_clk,
          mosi                        => pc_spi_mosi_out,
          miso                        => pc_spi_miso_in,
          cs_n                        => pc_spi_cs_out
        ) ;


      pc_flash_clk            <= '0' ;
      pc_flash_cs_out         <= '1' ;
      pc_flash_data_io        <= (others => '0') ;
      pc_flash_dir_out        <= '1' ;

    end generate use_PC ;

  no_use_PC:
    if (Collar_Control_usePC_c = '0') generate

      pc_spi_clk              <= '0' ;
      pc_spi_cs_out           <= '1' ;
      pc_spi_mosi_out         <= '0' ;

      pc_flash_clk            <= '0' ;
      pc_flash_cs_out         <= '1' ;
      pc_flash_data_io        <= (others => '0') ;
      pc_flash_dir_out        <= '1' ;

      StatCtlActive           <= '0' ;

    end generate no_use_PC ;

  --------------------------------------------------------------------------
  --  Event logging.
  --------------------------------------------------------------------------

  use_EventLogging:
    if (Collar_Control_useEventLogging_c = '1') generate

      component LoggingCounterArray is
        Generic (
          clk_freq_g            : natural     := 10e6 ;
          counter_size_g        : natural     := 8 ;
          address_size_g        : natural     := 9 ;
          counters_g            : natural     := 1 ;
          rollover_g            : std_logic   := '0'
        ) ;
        Port (
          reset                 : in    std_logic ;
          clk                   : in    std_logic ;
          mem_datafrom_in       : in    unsigned (counter_size_g-1 downto 0) ;
          mem_datato_out        : out   unsigned (counter_size_g-1 downto 0) ;
          mem_address_out       : out   unsigned (address_size_g-1 downto 0) ;
          mem_read_en_out       : out   std_logic ;
          mem_write_en_out      : out   std_logic ;
          counter_incr_in       : in    std_logic_vector (counters_g-1 downto 0) ;
          counter_clear_in      : in    std_logic ;
          counter_lock_in       : in    std_logic ;
          counters_changed_out  : out   std_logic ;
          busy_out              : out   std_logic
        ) ;
      end component LoggingCounterArray ;

      component eventmem IS
        PORT
        (
          address_a   : IN STD_LOGIC_VECTOR (eventcnt_addrbits_c-1 DOWNTO 0);
          address_b   : IN STD_LOGIC_VECTOR (eventcnt_addrbits_c-1 DOWNTO 0);
          clock_a     : IN STD_LOGIC  := '1';
          clock_b     : IN STD_LOGIC ;
          data_a      : IN STD_LOGIC_VECTOR (eventcnt_databits_c-1 DOWNTO 0);
          data_b      : IN STD_LOGIC_VECTOR (eventcnt_databits_c-1 DOWNTO 0);
          rden_a      : IN STD_LOGIC  := '1';
          rden_b      : IN STD_LOGIC  := '1';
          wren_a      : IN STD_LOGIC  := '0';
          wren_b      : IN STD_LOGIC  := '0';
          q_a         : OUT STD_LOGIC_VECTOR (eventcnt_databits_c-1 DOWNTO 0);
          q_b         : OUT STD_LOGIC_VECTOR (eventcnt_databits_c-1 DOWNTO 0)
        ) ;
      END component eventmem ;

      --  Constants and signals used to map to memory.

      signal evmemsrc_clk         : std_logic ;
      signal evmemsrc_readfrom    : std_logic_vector (eventcnt_databits_c-1
                                                      downto 0) ;
      signal evmemsrc_writeto     : std_logic_vector (eventcnt_databits_c-1
                                                      downto 0) ;
      signal evmemsrc_addr        : std_logic_vector (eventcnt_addrbits_c-1
                                                      downto 0) ;
      signal evmemsrc_read_en     : std_logic ;
      signal evmemsrc_write_en    : std_logic ;

    begin

      eventcnt : LoggingCounterArray
        Generic Map (
          clk_freq_g            => master_clk_freq_c,
          counter_size_g        => eventcnt_databits_c,
          address_size_g        => eventcnt_addrbits_c,
          counters_g            => eventcnt_events_c,
          rollover_g            => '0'
        )
        Port Map (
          reset                 => reset,
          clk                   => master_gated_clk,
          mem_datafrom_in       => unsigned (evmemsrc_readfrom),
          std_logic_vector (mem_datato_out)   => evmemsrc_writeto,
          std_logic_vector (mem_address_out)  => evmemsrc_addr,
          mem_read_en_out       => evmemsrc_read_en,
          mem_write_en_out      => evmemsrc_write_en,
          counter_incr_in       => eventcnt_incr,
          counter_clear_in      => eventcnt_clear,
          counter_lock_in       => eventcnt_lock,
          counters_changed_out  => eventcnt_changed,
          busy_out              => eventcnt_busy
        ) ;

      eventmemory : eventmem
        Port Map (
          address_a               => evmemsrc_addr,
          address_b               => evmemdst_addr,
          clock_a                 => master_gated_inv_clk,
          clock_b                 => evmemdst_clk,
          data_a                  => evmemsrc_writeto,
          data_b                  => evmemdst_writeto,
          rden_a                  => evmemsrc_read_en,
          rden_b                  => evmemdst_read_en,
          wren_a                  => evmemsrc_write_en,
          wren_b                  => evmemdst_write_en,
          q_a                     => evmemsrc_readfrom,
          q_b                     => evmemdst_readfrom
        ) ;

      --  Events mapping to the vector.

      ev_MainPowerSwitchOn        <=     CTL_MainPowerSwitch ;
      ev_MainPowerSwitchOff       <= not CTL_MainPowerSwitch ;
      ev_RechargeSwitchOn         <=     CTL_RechargeSwitch ;
      ev_RechargeSwitchOff        <= not CTL_RechargeSwitch ;
      ev_SolarCtlShutdownOn       <=     CTL_SolarCtlShutdown ;
      ev_SolarCtlShutdownOff      <= not CTL_SolarCtlShutdown ;
      ev_LevelShifter3p3On        <=     CTL_LevelShifter3p3 ;
      ev_LevelShifter3p3Off       <= not CTL_LevelShifter3p3 ;
      ev_LevelShifter1p8On        <=     CTL_LevelShifter1p8 ;
      ev_LevelShifter1p8Off       <= not CTL_LevelShifter1p8 ;
      ev_InertialOn1p8            <=     CTL_InertialOn1p8 ;
      ev_InertialOff2p5           <= not CTL_InertialOn2p5 ;
      ev_MicLeftOn                <=     CTL_MicLeftOn ;
      ev_MicLeftOff               <= not CTL_MicLeftOn ;
      ev_MicRightOn               <=     CTL_MicRightOn ;
      ev_MicRightOff              <= not CTL_MicRightOn ;
      ev_SDRAM_On                 <=     CTL_SDRAM_On ;
      ev_SDRAM_Off                <= not CTL_SDRAM_On ;
      ev_SDCardOn                 <=     CTL_SDCardOn ;
      ev_SDCardOff                <= not CTL_SDCardOn ;
      ev_GPS_On                   <=     CTL_GPS_On ;
      ev_GPS_Off                  <= not CTL_GPS_On ;
      ev_DataTX_On                <=     CTL_DataTX_On ;
      ev_DataTX_Off               <= not CTL_DataTX_On ;

      ev_BatteryGoodOn            <=     STAT_BatteryGood ;
      ev_BatteryGoodOff           <= not STAT_BatteryGood ;
      ev_SolarCtlOn               <=     STAT_SolarCtlOn ;
      ev_SolarCtlOff              <= not STAT_SolarCtlOn ;
      ev_BattMonLowOn             <=     STAT_BattMonLow ;
      ev_BattMonLowOff            <= not STAT_BattMonLow ;
      ev_ForceStartupOn           <=     STAT_ForceStartup ;
      ev_ForceStartupOff          <= not STAT_ForceStartup ;
      ev_PwrGood2p5On             <=     STAT_PwrGood2p5 ;
      ev_PwrGood2p5Off            <= not STAT_PwrGood2p5 ;
      ev_PwrGood3p3On             <=     STAT_PwrGood3p3 ;
      ev_PwrGood3p3Off            <= not STAT_PwrGood3p3 ;

    end generate use_EventLogging ;

  no_use_EventLogging:
    if (Collar_Control_useEventLogging_c = '0') generate

      eventcnt_changed      <= '0' ;
      eventcnt_busy         <= '0' ;
      evmemdst_readfrom     <= (others => '0') ;

    end generate no_use_EventLogging ;

  --------------------------------------------------------------------------
  --  SDRAM.
  --------------------------------------------------------------------------

  use_SDRAM:
    if (Collar_Control_useSDRAM_c = '1') generate

      --  Constants and signals used to map to memory buffers.

      constant inmem_rdwidth_c      : natural := 16 ;
      constant inmem_rdelements_c   : natural :=
                  8 * inmem_bytecnt_c / inmem_rdwidth_c ;
      constant inmem_rdaddrbits_c   : natural :=
                  const_bits (inmem_rdelements_c - 1) ;

      constant outmem_wrwidth_c     : natural := 16 ;
      constant outmem_wrelements_c  : natural :=
                  8 * outmem_bytecnt_c / outmem_wrwidth_c ;
      constant outmem_wraddrbits_c  : natural :=
                  const_bits (outmem_wrelements_c - 1) ;

      signal sdram_inrd_data  : std_logic_vector (inmem_rdwidth_c-1
                                                  downto 0) ;
      signal sdram_inrd_addr  : std_logic_vector (inmem_rdaddrbits_c-1
                                                  downto 0) ;
      signal sdram_inrd_en    : std_logic ;
      signal sdram_inrd_clk   : std_logic ;

      signal sdram_outwr_data : std_logic_vector (outmem_wrwidth_c-1
                                                  downto 0) ;
      signal sdram_outwr_addr : std_logic_vector (outmem_wraddrbits_c-1
                                                  downto 0) ;
      signal sdram_outwr_en   : std_logic ;
      signal sdram_outwr_clk  : std_logic ;

      --  Component declarations.

      component SDRAM_Controller is
        Generic (
          sysclk_freq_g         : natural     := 10e6 ;

          outmem_buffrows_g     : natural     := 1 ;
          outmem_buffcount_g    : natural     := 2 ;
          inmem_buffouts_g      : natural     := 1 ;
          inmem_buffcount_g     : natural     := 2 ;
          sdram_space_g         : SDRAM_Capacity_t  := SDRAM_32_Capacity_c ;
          sdram_times_g         : SDRAM_Timing_t    := SDRAM_75_3_Timing_c
        ) ;
        Port (
          reset                 : in    std_logic ;
          sysclk                : in    std_logic ;

          ready_out             : out   std_logic ;

          inmem_buffready_in    : in    std_logic ;
          inmem_datafrom_in     : in    std_logic_vector (sdram_space_g.DATABITS-1
                                                          downto 0) ;
          inmem_address_out     : out
              std_logic_vector (const_bits (inmem_buffcount_g * inmem_buffouts_g *
                                            outmem_buffrows_g *
                                            sdram_space_g.ROWBITS /
                                            sdram_space_g.DATABITS - 1) - 1
                                              downto 0) ;
          inmem_read_en_out     : out   std_logic ;
          inmem_clk_out         : out   std_logic ;

          outmem_buffready_in   : in    std_logic ;
          outmem_datato_out     : out   std_logic_vector (sdram_space_g.DATABITS-1
                                                          downto 0) ;
          outmem_address_out    : out
              std_logic_vector (const_bits (outmem_buffcount_g *
                                            outmem_buffrows_g *
                                            sdram_space_g.ROWBITS /
                                            sdram_space_g.DATABITS - 1) - 1
                                              downto 0) ;
          outmem_write_en_out   : out   std_logic ;
          outmem_clk_out        : out   std_logic ;
          outmem_amt_out        : out
              unsigned (const_bits (sdram_space_g.BANKS * sdram_space_g.ROWCOUNT *
                                    sdram_space_g.ROWBITS / 8 - 1) - 1 downto 0) ;
          outmem_writing_out    : out   std_logic ;

          sdram_data_in         : in    std_logic_vector (sdram_space_g.DATABITS-1
                                                            downto 0) ;
          sdram_data_out        : out   std_logic_vector (sdram_space_g.DATABITS-1
                                                            downto 0) ;
          sdram_data_dir        : out   std_logic ;

          sdram_mask_out        : out
              std_logic_vector (sdram_space_g.DATABITS / 8 - 1 downto 0) ;
          sdram_address_out     : out   unsigned (sdram_space_g.ADDRBITS-1
                                                            downto 0) ;
          sdram_bank_out        : out
              unsigned (const_bits (sdram_space_g.BANKS - 1)-1 downto 0) ;
          sdram_command_out     : out   std_logic_vector (sdram_space_g.CMDBITS-1
                                                            downto 0) ;
          sdram_clk_en_out      : out   std_logic ;
          sdram_clk_out         : out   std_logic ;
          sdram_empty_out       : out   std_logic ;
          sdram_forceout_in     : in    std_logic
        ) ;
      end component SDRAM_Controller ;

      component outmem IS
        PORT
        (
          data        : IN STD_LOGIC_VECTOR (outmem_wrwidth_c-1 DOWNTO 0) ;
          rdaddress   : IN STD_LOGIC_VECTOR (outmem_rdaddrbits_c-1 DOWNTO 0) ;
          rdclock     : IN STD_LOGIC ;
          rden        : IN STD_LOGIC  := '1' ;
          wraddress   : IN STD_LOGIC_VECTOR (outmem_wraddrbits_c-1 DOWNTO 0) ;
          wrclock     : IN STD_LOGIC  := '1' ;
          wren        : IN STD_LOGIC  := '0' ;
          q           : OUT STD_LOGIC_VECTOR (outmem_rdwidth_c-1 DOWNTO 0)
        ) ;
      END component outmem ;

      component inmem IS
        PORT
        (
          data        : IN STD_LOGIC_VECTOR (inmem_wrwidth_c-1 DOWNTO 0) ;
          rdaddress   : IN STD_LOGIC_VECTOR (inmem_rdaddrbits_c-1 DOWNTO 0) ;
          rdclock     : IN STD_LOGIC ;
          rden        : IN STD_LOGIC  := '1' ;
          wraddress   : IN STD_LOGIC_VECTOR (inmem_wraddrbits_c-1 DOWNTO 0) ;
          wrclock     : IN STD_LOGIC  := '1' ;
          wren        : IN STD_LOGIC  := '0' ;
          q           : OUT STD_LOGIC_VECTOR (inmem_rdwidth_c-1 DOWNTO 0)
        ) ;
      END component inmem ;

      --  Signals used for mapping to the device.

      signal sdram_clock      : std_logic ;
      signal sdram_clk_en     : std_logic ;
      signal sdram_command    : std_logic_vector (sdram_command_out'length-1
                                                  downto 0) ;
      signal sdram_mask       : std_logic_vector (sdram_mask_out'length-1
                                                  downto 0) ;
      signal sdram_bank       : std_logic_vector (sdram_bank_out'length-1
                                                  downto 0) ;
      signal sdram_addr       : std_logic_vector (sdram_addr_out'length-1
                                                  downto 0) ;
      signal sdram_indata     : std_logic_vector (sdram_data_io'length-1
                                                  downto 0) ;
      signal sdram_outdata    : std_logic_vector (sdram_data_io'length-1
                                                  downto 0) ;
      signal sdram_dirdata    : std_logic ;

    begin

      sdcard_buffer : SDRAM_Controller
        Generic Map (
          sysclk_freq_g         => master_clk_freq_c,

          outmem_buffrows_g     => outmem_buffrows_c,
          outmem_buffcount_g    => outmem_buffcount_c,
          inmem_buffouts_g      => inmem_buffouts_c,
          inmem_buffcount_g     => inmem_buffcount_c,
          sdram_space_g         => sdram_space_g,
          sdram_times_g         => sdram_times_g
        )
        Port Map (
          reset                 => reset or not CTL_SDRAM_On,
          sysclk                => master_clk,
          ready_out             => sdram_ready,

          inmem_buffready_in    => sdram_inready,
          inmem_datafrom_in     => sdram_inrd_data,
          inmem_address_out     => sdram_inrd_addr,
          inmem_read_en_out     => sdram_inrd_en,
          inmem_clk_out         => sdram_inrd_clk,

          outmem_buffready_in   => sdram_outready,
          outmem_datato_out     => sdram_outwr_data,
          outmem_address_out    => sdram_outwr_addr,
          outmem_write_en_out   => sdram_outwr_en,
          outmem_clk_out        => sdram_outwr_clk,
          outmem_amt_out        => sdram_outamt,
          outmem_writing_out    => sdram_outwriting,

          sdram_data_in         => sdram_indata,
          sdram_data_out        => sdram_outdata,
          sdram_data_dir        => sdram_dirdata,

          sdram_mask_out        => sdram_mask,
          std_logic_vector (sdram_address_out)  => sdram_addr,
          std_logic_vector (sdram_bank_out)     => sdram_bank,
          sdram_command_out     => sdram_command,
          sdram_clk_en_out      => sdram_clk_en,
          sdram_clk_out         => sdram_clock,
          sdram_empty_out       => sdram_empty,
          sdram_forceout_in     => sdram_forceout
        ) ;

      sdcard_buffout : outmem
        Port Map (
          data        => sdram_outwr_data,
          rdaddress   => sdram_outrd_addr,
          rdclock     => sdram_outrd_clk,
          rden        => sdram_outrd_en,
          wraddress   => sdram_outwr_addr,
          wrclock     => sdram_outwr_clk,
          wren        => sdram_outwr_en,
          q           => sdram_outrd_data
        ) ;

      sdcard_buffin : inmem
        Port Map (
          data        => sdram_inwr_data,
          rdaddress   => sdram_inrd_addr,
          rdclock     => sdram_inrd_clk,
          rden        => sdram_inrd_en,
          wraddress   => sdram_inwr_addr,
          wrclock     => sdram_inwr_clk,
          wren        => sdram_inwr_en,
          q           => sdram_inrd_data
        ) ;

      ----------------------------------------------------------------------
      --  All I/O lines forced low when device is off, otherwise they are
      --  driven from the component.
      ----------------------------------------------------------------------

      sdram_indata            <= sdram_data_io ;

      sdram_on : process (CTL_SDRAM_On, sdram_clock, sdram_clk_en,
                          sdram_command, sdram_mask, sdram_bank,
                          sdram_addr, sdram_outdata, sdram_dirdata)
      begin
        if (CTL_SDRAM_On = '0') then
          sdram_clk           <= '0' ;
          sdram_clk_en_out    <= '0' ;
          sdram_command_out   <= (others => '0') ;
          sdram_mask_out      <= (others => '0') ;
          sdram_bank_out      <= (others => '0') ;
          sdram_addr_out      <= (others => '0') ;
          sdram_data_io       <= (others => '0') ;
        else
          sdram_clk           <= sdram_clock ;
          sdram_clk_en_out    <= sdram_clk_en ;
          sdram_command_out   <= sdram_command ;
          sdram_mask_out      <= sdram_mask ;
          sdram_bank_out      <= sdram_bank ;
          sdram_addr_out      <= sdram_addr ;

          if (sdram_dirdata = '1') then
            sdram_data_io     <= sdram_outdata ;
          else
            sdram_data_io     <= (others => 'Z') ;
          end if ;
        end if ;
      end process sdram_on ;

  end generate use_SDRAM ;

  no_use_SDRAM:
    if (Collar_Control_useSDRAM_c = '0') generate

      sdram_clk               <= '0' ;
      sdram_clk_en_out        <= '0' ;
      sdram_command_out       <= (others => '0') ;
      sdram_mask_out          <= (others => '0') ;
      sdram_bank_out          <= (others => '0') ;
      sdram_addr_out          <= (others => '0') ;
      sdram_data_io           <= (others => '0') ;

      sdram_ready             <= '1' ;
      sdram_empty             <= '0' ;

      sdram_outwriting        <= '0' ;
      sdram_outamt            <= (others => '0') ;
      sdram_outrd_data        <= (others => '0') ;

    end generate no_use_SDRAM ;

  --------------------------------------------------------------------------
  --  SD Card controller.
  --------------------------------------------------------------------------

  use_SD:
    if (Collar_Control_useSD_c = '1') generate

      component microsd_controller_dir is
        generic(

          clk_freq_g                :natural    := 50E6;
          buf_size_g                :natural    := 2048;
          block_size_g              :natural    := 512;
          hs_sdr25_mode_g            :std_logic  := '1';
          clk_divide_g              :natural    := 128;
          signalling_18_en_g        :std_logic  := '0'
        );

        port(

          rst_n           :in      std_logic;
          clk             :in      std_logic;
          clock_enable    :in      std_logic;
          data_input      :in      std_logic_vector(7 downto 0);
          data_we         :in      std_logic;
          data_full       :out     std_logic;
          data_sd_start_address     :in      std_logic_vector(31 downto 0);
          data_nblocks              :in      std_logic_vector(31 downto 0);

          data_current_block_written      :out     std_logic_vector(31 downto 0);
          sd_block_written_flag           :out     std_logic;
          buffer_level                    :out     std_logic_vector (natural(trunc(log2(
                                          real(buf_size_g/block_size_g)))) downto 0);

          sd_clk                          :out     std_logic;

          sd_cmd_in                       : in      std_logic ;
          sd_cmd_out                      : out     std_logic ;
          sd_cmd_dir                      : out     std_logic ;
          sd_dat_in                       : in      std_logic_vector (3 downto 0) ;
          sd_dat_out                      : out     std_logic_vector (3 downto 0) ;
          sd_dat_dir                      : out     std_logic_vector (3 downto 0) ;

          v_3_3_on_off                    :out     std_logic;
          v_1_8_on_off                    :out     std_logic;

          init_start                      :in     std_logic;
          user_led_n_out                  :out    std_logic_vector(3 downto 0);
          ext_trigger                     :out    std_logic

        );
      end component microsd_controller_dir ;

    component sd_loader is
      generic(
        OUTMEM_BUFFROWS       : natural     := 1 ;
        OUTMEM_BUFFCOUNT      : natural     := 2 ;
        sdram_space_g         : SDRAM_Capacity_t  := SDRAM_16_Capacity_c;
        sdram_outbuf_size_bytes_g : natural := 4096;
        buf_size_g            :   natural := 2048;
        block_size_g          :   natural := 512;
        enable_magmem_g       :   std_logic := '0'
      );
      port(

        clk        : in std_logic;
        rst_n      : in std_logic;

        startup_in              : in std_logic;

        data_nbytes_in          : in std_logic_vector (const_bits (sdram_space_g.BANKS * sdram_space_g.ROWCOUNT *
                                sdram_space_g.ROWBITS / 8 - 1) - 1 downto 0) ;
        outbuf_data_rdy_in      : in std_logic;

        outbuf_sd_q_b_in        : in std_logic_vector(7 downto 0);
        sd_outbuf_rd_en_b_out   : out std_logic;
        sd_outbuf_clk_b_out     : out std_logic;
        sd_outbuf_address_b_out : out std_logic_vector(natural(trunc(log2(real(sdram_outbuf_size_bytes_g-1)))) downto 0);

        sd_outmem_buffready_out : out std_logic;

        mem_req_a_out           : out std_logic;
        mem_rec_a_in            : in std_logic;


        sd_magram_clk_a_out     : out std_logic;
        sd_magram_wr_en_a_out   : out std_logic;
        sd_magram_rd_en_a_out   : out std_logic;
        sd_magram_address_a_out : out std_logic_vector(natural(trunc(log2(real(
                                (magmem_buffer_bytes/magmem_buffer_num)-1)))) downto 0);
        sd_magram_data_a_out    : out std_logic_vector(7 downto 0);
        magram_sd_q_a_in        : in std_logic_vector(7 downto 0);

        dw_en                   : in std_logic;
        crit_block_serviced     : out std_logic;

        data_input                         :out      std_logic_vector(7 downto 0);
        data_we                            :out      std_logic;
        data_full                          :in       std_logic;
        data_sd_start_address              :out      std_logic_vector(31 downto 0);
        data_nblocks                       :out      std_logic_vector(31 downto 0);
        data_current_block_written         :in       std_logic_vector(31 downto 0);
        sd_block_written_flag              :in       std_logic;
        buffer_level                       :in       std_logic_vector (natural(trunc(log2(real(buf_size_g/block_size_g)))) downto 0);

        blocks_past_crit                   :in std_logic_vector(7 downto 0)

      );
    end component;

      --  SD loader to Magnetic Memory communications signals.

      signal sdl_magmem_clk       : std_logic ;
      signal sdl_magmem_wr_en     : std_logic ;
      signal sdl_magmem_rd_en     : std_logic ;
       signal sdl_magmem_addr      : std_logic_vector(natural(trunc(log2(real((magmem_buffer_bytes/magmem_buffer_num)-1)))) downto 0);
      --signal sdl_magmem_addr      : std_logic_vector (magmem_addrbits_c-1
      --                                                downto 0) ;
      signal sdl_magmem_writeto   : std_logic_vector (magmem_databits_c-1
                                                      downto 0) ;
      signal sdl_magmem_control   : std_logic_vector (magmem_iobits_c-1
                                                      downto 0) ;

      --  SD loader to SD Card controller communication signals.

      constant outmem_buffblks_c  : natural := sdram_rowbytes_c /
                                               sdcard_blksize_c ;

      signal sdl_sdcard_writeto   : std_logic_vector (7 downto 0) ;
      signal sdl_sdcard_wr_en     : std_logic ;
      signal sdl_sdcard_full      : std_logic ;
      signal sdl_sdcard_startblk  : std_logic_vector (sdcard_blknobits_c-1
                                                      downto 0) ;
      signal sdl_sdcard_nblocks   : std_logic_vector (sdcard_blknobits_c-1
                                                      downto 0) ;
      signal sdl_sdcard_lastblk   : std_logic_vector (sdcard_blknobits_c-1
                                                      downto 0) ;
      signal sdl_sdcard_lastflag  : std_logic ;
      signal sdl_sdcard_bufflevel :
                std_logic_vector (const_bits (outmem_buffblks_c-1)
                                  downto 0) ;
      signal sdl_sdcard_critdone  : std_logic ;
      signal sdl_sdcard_critpast  : std_logic_vector (7 downto 0) ;

      --  Signals for I/O mapping.

      signal sd_clock     : std_logic ;
      signal sd_incmd     : std_logic ;
      signal sd_outcmd    : std_logic ;
      signal sd_dircmd    : std_logic ;
      signal sd_indata    : std_logic_vector (sd_data_io'length-1
                                              downto 0) ;
      signal sd_outdata   : std_logic_vector (sd_data_io'length-1
                                              downto 0) ;
      signal sd_dirdata   : std_logic_vector (sd_data_io'length-1
                                              downto 0) ;

    begin

      --  SD Card Loader mapping.

      sdload : sd_loader
        generic map (
          OUTMEM_BUFFROWS           => outmem_buffrows_c,
          OUTMEM_BUFFCOUNT          => outmem_buffcount_c,
          sdram_space_g               => sdram_space_g,
          sdram_outbuf_size_bytes_g => outmem_bytecnt_c,
          buf_size_g                => sdram_rowbytes_c,
          block_size_g              => sdcard_blksize_c
        )
        port map (
          clk                       => master_clk,
          rst_n                     => (not reset) and CTL_SDCardOn,
          startup_in                => sdcard_start,
          data_nbytes_in            => std_logic_vector (sdram_outamt),
          outbuf_data_rdy_in        => sdram_outwriting,
          outbuf_sd_q_b_in          => sdram_outrd_data,
          sd_outbuf_rd_en_b_out     => sdram_outrd_en,
          sd_outbuf_clk_b_out       => sdram_outrd_clk,
          sd_outbuf_address_b_out   => sdram_outrd_addr,
          sd_outmem_buffready_out   => sdram_outready,
          mem_req_a_out             => magmem_requesters (magmemrq_sdcard_c),
          mem_rec_a_in              => magmem_receivers  (magmemrq_sdcard_c),
          sd_magram_clk_a_out       => sdl_magmem_clk,
          sd_magram_wr_en_a_out     => sdl_magmem_wr_en,
          sd_magram_rd_en_a_out     => sdl_magmem_rd_en,
          sd_magram_address_a_out   => sdl_magmem_addr,
          sd_magram_data_a_out      => sdl_magmem_writeto,
          magram_sd_q_a_in          => magmemsrc_readfrom,
          data_input                => sdl_sdcard_writeto,
          data_we                   => sdl_sdcard_wr_en,
          data_full                 => sdl_sdcard_full,
          data_sd_start_address     => sdl_sdcard_startblk,
          data_nblocks              => sdl_sdcard_nblocks,
          data_current_block_written  => sdl_sdcard_lastblk,
          sd_block_written_flag     => sdl_sdcard_lastflag,
          buffer_level              => sdl_sdcard_bufflevel,
          dw_en                     => '0',
          crit_block_serviced       => sdl_sdcard_critdone,
          blocks_past_crit          => sdl_sdcard_critpast
        );



      sdl_magmem_control    <= master_gated_inv_clk &
                               sdl_magmem_wr_en     & sdl_magmem_rd_en &
                               sdl_magmem_writeto   & mm_buffno &
                               sdl_magmem_addr ;

      set2D_element (magmemrq_sdcard_c, sdl_magmem_control,
                     magmem_input_tbl) ;

      --  SD Card mapping.

      sdcard : microsd_controller_dir
        generic map (
          clk_freq_g          => master_clk_freq_c,
          buf_size_g        => sdcard_blksize_c * 4,
          block_size_g      => sdcard_blksize_c,
          hs_sdr25_mode_g     => '1',
          clk_divide_g        => natural (real (master_clk_freq_c) / 400000.0)
        )
        port map (
          rst_n                       => (not reset) and CTL_SDCardOn,
          clk                         => master_clk,
          clock_enable                => '1',

          data_input                  => sdl_sdcard_writeto,
          data_we                     => sdl_sdcard_wr_en,
          data_full                   => sdl_sdcard_full,
          data_sd_start_address       => sdl_sdcard_startblk,
          data_nblocks                => sdl_sdcard_nblocks,
          data_current_block_written  => sdl_sdcard_lastblk,
          sd_block_written_flag       => sdl_sdcard_lastflag,

          sd_clk                      => sd_clk,
          sd_cmd_in                   => sd_incmd,
          sd_cmd_out                  => sd_outcmd,
          sd_cmd_dir                  => sd_dircmd,
          sd_dat_in                   => sd_indata,
          sd_dat_out                  => sd_outdata,
          sd_dat_dir                  => sd_dirdata,

          V_3_3_ON_OFF                => CTL_LevelShifter3p3,
          V_1_8_ON_OFF                => CTL_LevelShifter1p8,

          init_start                  => not sdcard_start
        ) ;

      ----------------------------------------------------------------------
      --  All I/O lines forced low when device is off, otherwise they are
      --  driven from the component.
      ----------------------------------------------------------------------

      sd_incmd                <= sd_cmd_io ;
      sd_indata               <= sd_data_io ;

      sdcard_on : process (CTL_SDCardOn, sd_clock,
                           sd_dircmd,  sd_outcmd,
                           sd_dirdata, sd_outdata)
      begin
        if (CTL_SDCardOn = '0') then
          sd_clk              <= '0' ;
          sd_cmd_io           <= '0' ;
          sd_data_io          <= (others => '0') ;
        else
          sd_clk              <= sd_clock ;

          if (sd_dircmd = '1') then
            sd_cmd_io         <= sd_outcmd ;
          else
            sd_cmd_io         <= 'Z' ;
          end if ;

          for i in 0 to sd_dirdata'length-1 loop
            if (sd_dirdata (i) = '1') then
              sd_data_io (i)  <= sd_outdata (i) ;
            else
              sd_data_io (i)  <= 'Z' ;
            end if ;
          end loop ;
        end if ;
      end process sdcard_on ;

    end generate use_SD ;

  no_use_SD:
    if (Collar_Control_useSD_c = '0') generate

      sd_clk        <= '0' ;
      sd_cmd_io     <= '0' ;
      sd_data_io    <= (others => '0') ;

    end generate no_use_SD ;

  --------------------------------------------------------------------------
  --  Direct connect SD Card controller.  Does not use voltage level
  --  shifting.
  --------------------------------------------------------------------------

  use_SDH:
    if (Collar_Control_useSDH_c = '1') generate

      component microsd_controller_dir is
        generic(

          clk_freq_g                :natural    := 50E6;
          buf_size_g                :natural    := 2048;
          block_size_g              :natural    := 512;
          hs_sdr25_mode_g            :std_logic  := '1';
          clk_divide_g              :natural    := 128;
          signalling_18_en_g        :std_logic  := '0'
        );

        port(

          rst_n           :in      std_logic;
          clk             :in      std_logic;
          clock_enable    :in      std_logic;
          data_input      :in      std_logic_vector(7 downto 0);
          data_we         :in      std_logic;
          data_full       :out     std_logic;
          data_sd_start_address     :in      std_logic_vector(31 downto 0);
          data_nblocks              :in      std_logic_vector(31 downto 0);

          data_current_block_written      :out     std_logic_vector(31 downto 0);
          sd_block_written_flag           :out     std_logic;
          buffer_level                    :out     std_logic_vector (natural(trunc(log2(
                                          real(buf_size_g/block_size_g)))) downto 0);

          sd_clk                          :out     std_logic;

          sd_cmd_in                       : in      std_logic ;
          sd_cmd_out                      : out     std_logic ;
          sd_cmd_dir                      : out     std_logic ;
          sd_dat_in                       : in      std_logic_vector (3 downto 0) ;
          sd_dat_out                      : out     std_logic_vector (3 downto 0) ;
          sd_dat_dir                      : out     std_logic_vector (3 downto 0) ;

          v_3_3_on_off                    :out     std_logic;
          v_1_8_on_off                    :out     std_logic;

          init_start                      :in     std_logic;
          user_led_n_out                  :out    std_logic_vector(3 downto 0);
          ext_trigger                     :out    std_logic

        );
      end component microsd_controller_dir ;

      -- component sd_loader is
        -- generic (
          -- OUTMEM_BUFFROWS       : natural     := 1 ;
          -- OUTMEM_BUFFCOUNT      : natural     := 2 ;
          -- SDRAM_SPACE           : SDRAM_Capacity_t  := SDRAM_32_Capacity_c;
          -- sdram_outbuf_size_bytes_g : natural := 4096;
          -- buf_size_g            :   natural := 2048;
          -- block_size_g          :   natural := 512
        -- );
        -- port (
          -- clk        : in std_logic;
          -- rst_n      : in std_logic;
          -- startup_in              : in std_logic;
          -- data_nbytes_in          : in std_logic_vector(const_bits (SDRAM_SPACE.BANKS * SDRAM_SPACE.ROWCOUNT *
                                    -- SDRAM_SPACE.ROWBITS / 8 - 1) - 1 downto 0) ;
          -- outbuf_data_rdy_in      : in std_logic;
          -- outbuf_sd_q_b_in        : in std_logic_vector(7 downto 0);
          -- sd_outbuf_rd_en_b_out   : out std_logic;
          -- sd_outbuf_address_b_out : out std_logic_vector(natural(trunc(log2(real(sdram_outbuf_size_bytes_g-1)))) downto 0);
          -- mem_req_a_out           : out std_logic;
          -- mem_rec_a_in            : in std_logic;
          -- sd_magram_wr_en_a_out   : out std_logic;
          -- sd_magram_rd_en_a_out   : out std_logic;
          -- sd_magram_address_a_out : out std_logic_vector(natural(trunc(log2(real(magmem_buffer_bytes-1)))) downto 0);
          -- sd_magram_data_a_out    : out std_logic_vector(7 downto 0);
          -- magram_sd_q_a_in        : in std_logic_vector(7 downto 0);
          -- dw_en                   : in std_logic;
          -- crit_block_serviced     : out std_logic;
          -- data_input                         :out      std_logic_vector(7 downto 0);
          -- data_we                            :out      std_logic;
          -- data_full                          :in       std_logic;
          -- data_sd_start_address              :out      std_logic_vector(31 downto 0);
          -- data_nblocks                       :out      std_logic_vector(31 downto 0);
          -- data_current_block_written         :in       std_logic_vector(31 downto 0);
          -- sd_block_written_flag              :in       std_logic;
          -- buffer_level                       :in       std_logic_vector (natural(trunc(log2(real(buf_size_g/block_size_g)))) downto 0);
          -- blocks_past_crit                   :in std_logic_vector(7 downto 0)
        -- );
      -- end component sd_loader;

    component sd_loader is
      generic(
        OUTMEM_BUFFROWS       : natural     := 1 ;
        OUTMEM_BUFFCOUNT      : natural     := 2 ;
        sdram_space_g         : SDRAM_Capacity_t  := SDRAM_16_Capacity_c;
        sdram_outbuf_size_bytes_g : natural := 4096;
        buf_size_g            :   natural := 2048;
        block_size_g          :   natural := 512;
        enable_magmem_g       :   std_logic := '0'
      );
      port(

        clk        : in std_logic;
        rst_n      : in std_logic;

        startup_in              : in std_logic;

        data_nbytes_in          : in std_logic_vector (const_bits (sdram_space_g.BANKS * sdram_space_g.ROWCOUNT *
                                sdram_space_g.ROWBITS / 8 - 1) - 1 downto 0) ;
        outbuf_data_rdy_in      : in std_logic;

        outbuf_sd_q_b_in        : in std_logic_vector(7 downto 0);
        sd_outbuf_rd_en_b_out   : out std_logic;
        sd_outbuf_clk_b_out     : out std_logic;
        sd_outbuf_address_b_out : out std_logic_vector(natural(trunc(log2(real(sdram_outbuf_size_bytes_g-1)))) downto 0);

        sd_outmem_buffready_out : out std_logic;

        mem_req_a_out           : out std_logic;
        mem_rec_a_in            : in std_logic;


        sd_magram_clk_a_out     : out std_logic;
        sd_magram_wr_en_a_out   : out std_logic;
        sd_magram_rd_en_a_out   : out std_logic;
        sd_magram_address_a_out : out std_logic_vector(natural(trunc(log2(
                                      real((magmem_buffer_bytes/magmem_buffer_num)-1)
                                      ))) downto 0);
        sd_magram_data_a_out    : out std_logic_vector(7 downto 0);
        magram_sd_q_a_in        : in std_logic_vector(7 downto 0);

        dw_en                   : in std_logic;
        crit_block_serviced     : out std_logic;

        data_input                         :out      std_logic_vector(7 downto 0);
        data_we                            :out      std_logic;
        data_full                          :in       std_logic;
        data_sd_start_address              :out      std_logic_vector(31 downto 0);
        data_nblocks                       :out      std_logic_vector(31 downto 0);
        data_current_block_written         :in       std_logic_vector(31 downto 0);
        sd_block_written_flag              :in       std_logic;
        buffer_level                       :in       std_logic_vector (natural(trunc(log2(real(buf_size_g/block_size_g)))) downto 0);

        blocks_past_crit                   :in std_logic_vector(7 downto 0)

      );
    end component;

      --  SD loader to Magnetic Memory communications signals.

      signal sdl_magmem_clk       : std_logic ;
      signal sdl_magmem_wr_en     : std_logic ;
      signal sdl_magmem_rd_en     : std_logic ;

      signal sdl_magmem_addr      : std_logic_vector(natural(trunc(log2(real((magmem_buffer_bytes/magmem_buffer_num)-1)))) downto 0);

      -- signal sdl_magmem_addr      : std_logic_vector (magmem_addrbits_c-1
                                                      -- downto 0) ;
      signal sdl_magmem_writeto   : std_logic_vector (magmem_databits_c-1
                                                      downto 0) ;
      signal sdl_magmem_control   : std_logic_vector (magmem_iobits_c-1
                                                      downto 0) ;

      --  SD loader to SD Card controller communication signals.

      constant outmem_buffblks_c  : natural := sdram_rowbytes_c /
                                               sdcard_blksize_c ;

      signal sdl_sdcard_writeto   : std_logic_vector (7 downto 0) ;
      signal sdl_sdcard_wr_en     : std_logic ;
      signal sdl_sdcard_full      : std_logic ;
      signal sdl_sdcard_startblk  : std_logic_vector (sdcard_blknobits_c-1
                                                      downto 0) ;
      signal sdl_sdcard_nblocks   : std_logic_vector (sdcard_blknobits_c-1
                                                      downto 0) ;
      signal sdl_sdcard_lastblk   : std_logic_vector (sdcard_blknobits_c-1
                                                      downto 0) ;
      signal sdl_sdcard_lastflag  : std_logic ;
      signal sdl_sdcard_bufflevel :
                std_logic_vector (const_bits (outmem_buffblks_c-1)
                                  downto 0) ;
      signal sdl_sdcard_critdone  : std_logic ;
      signal sdl_sdcard_critpast  : std_logic_vector (7 downto 0) ;

      --  Signals for I/O mapping.

      signal sd_clock     : std_logic ;
      signal sd_incmd     : std_logic ;
      signal sd_outcmd    : std_logic ;
      signal sd_dircmd    : std_logic ;
      signal sd_indata    : std_logic_vector (sd_data_io'length-1
                                              downto 0) ;
      signal sd_outdata   : std_logic_vector (sd_data_io'length-1
                                              downto 0) ;
      signal sd_dirdata   : std_logic_vector (sd_data_io'length-1
                                              downto 0) ;

    begin

      --  SD Card Loader mapping.

      sdload : sd_loader
        generic map (
          OUTMEM_BUFFROWS           => outmem_buffrows_c,
          OUTMEM_BUFFCOUNT          => outmem_buffcount_c,
          sdram_space_g               => sdram_space_g,
          sdram_outbuf_size_bytes_g => outmem_bytecnt_c,
          buf_size_g                => sdram_rowbytes_c,
          block_size_g              => sdcard_blksize_c
        )
        port map (
          clk                       => master_clk,
          rst_n                     => (not reset) and CTL_SDCardOn,
          startup_in                => sdcard_start,
          data_nbytes_in            => std_logic_vector (sdram_outamt),
          outbuf_data_rdy_in        => sdram_outwriting,
          outbuf_sd_q_b_in          => sdram_outrd_data,
          sd_outbuf_rd_en_b_out     => sdram_outrd_en,
          sd_outbuf_clk_b_out       => sdram_outrd_clk,
          sd_outbuf_address_b_out   => sdram_outrd_addr,
          sd_outmem_buffready_out   => sdram_outready,
          mem_req_a_out             => magmem_requesters (magmemrq_sdcard_c),
          mem_rec_a_in              => magmem_receivers  (magmemrq_sdcard_c),
          sd_magram_clk_a_out       => sdl_magmem_clk,
          sd_magram_wr_en_a_out     => sdl_magmem_wr_en,
          sd_magram_rd_en_a_out     => sdl_magmem_rd_en,
          sd_magram_address_a_out   => sdl_magmem_addr,
          sd_magram_data_a_out      => sdl_magmem_writeto,
          magram_sd_q_a_in          => magmemsrc_readfrom,
          data_input                => sdl_sdcard_writeto,
          data_we                   => sdl_sdcard_wr_en,
          data_full                 => sdl_sdcard_full,
          data_sd_start_address     => sdl_sdcard_startblk,
          data_nblocks              => sdl_sdcard_nblocks,
          data_current_block_written  => sdl_sdcard_lastblk,
          sd_block_written_flag     => sdl_sdcard_lastflag,
          buffer_level              => sdl_sdcard_bufflevel,
          dw_en                     => '0',
          crit_block_serviced       => sdl_sdcard_critdone,
          blocks_past_crit          => sdl_sdcard_critpast
        );

      sdl_magmem_control    <= master_gated_inv_clk &
                               sdl_magmem_wr_en     & sdl_magmem_rd_en &
                               sdl_magmem_writeto   & mm_buffno &
                               sdl_magmem_addr ;

      set2D_element (magmemrq_sdcard_c, sdl_magmem_control,
                     magmem_input_tbl) ;

      --  SD Card mapping.

      sdcard : microsd_controller_dir
        generic map (
          clk_freq_g          => master_clk_freq_c,
          buf_size_g        => sdcard_blksize_c * 4,
          block_size_g      => sdcard_blksize_c,
          hs_sdr25_mode_g     => '1',
          clk_divide_g        => natural (real (master_clk_freq_c) / 400000.0)
        )
        port map (
          rst_n                       => (not reset) and CTL_SDCardOn,
          clk                         => master_clk,
          clock_enable                => '1',

          data_input                  => sdl_sdcard_writeto,
          data_we                     => sdl_sdcard_wr_en,
          data_full                   => sdl_sdcard_full,
          data_sd_start_address       => sdl_sdcard_startblk,
          data_nblocks                => sdl_sdcard_nblocks,
          data_current_block_written  => sdl_sdcard_lastblk,
          sd_block_written_flag       => sdl_sdcard_lastflag,

          sd_clk                      => sd_clock,
          sd_cmd_in                   => sd_incmd,
          sd_cmd_out                  => sd_outcmd,
          sd_cmd_dir                  => sd_dircmd,
          sd_dat_in                   => sd_indata,
          sd_dat_out                  => sd_outdata,
          sd_dat_dir                  => sd_dirdata,

          init_start                  => not sdcard_start
        ) ;

      ----------------------------------------------------------------------
      --  All I/O lines forced low when device is off, otherwise they are
      --  driven from the component.
      ----------------------------------------------------------------------

      sd_incmd                <= sdh_cmd_io ;
      sd_indata               <= sdh_data_io ;

      sdcard_on : process (CTL_SDCardOn, sd_clock,
                           sd_dircmd,  sd_outcmd,
                           sd_dirdata, sd_outdata)
      begin
        if (CTL_SDCardOn = '0') then
          sdh_clk             <= '0' ;
          sdh_cmd_io          <= '0' ;
          sdh_data_io         <= (others => '0') ;
        else
          sdh_clk             <= sd_clock ;

          if (sd_dircmd = '1') then
            sdh_cmd_io        <= sd_outcmd ;
          else
            sdh_cmd_io        <= 'Z' ;
          end if ;

          for i in 0 to sd_dirdata'length-1 loop
            if (sd_dirdata (i) = '1') then
              sdh_data_io (i) <= sd_outdata (i) ;
            else
              sdh_data_io (i) <= 'Z' ;
            end if ;
          end loop ;
        end if ;
      end process sdcard_on ;

  end generate use_SDH ;

  no_use_SDH:
    if (Collar_Control_useSDH_c = '0') generate

      sdh_clk        <= '0' ;
      sdh_cmd_io     <= '0' ;
      sdh_data_io    <= (others => '0') ;

  end generate no_use_SDH ;

  --------------------------------------------------------------------------
  --  GPS RAM
  --------------------------------------------------------------------------

  use_GPS_RAM:
    if (Collar_Control_useGPSRAM_c = '1') generate

      component gps_ram IS
        PORT
        (
          address_a   : IN STD_LOGIC_VECTOR (gpsmem_addrbits_c-1 DOWNTO 0);
          address_b   : IN STD_LOGIC_VECTOR (gpsmem_addrbits_c-1 DOWNTO 0);
          clock_a     : IN STD_LOGIC  := '1';
          clock_b     : IN STD_LOGIC ;
          data_a      : IN STD_LOGIC_VECTOR (gpsmem_databits_c-1 DOWNTO 0);
          data_b      : IN STD_LOGIC_VECTOR (gpsmem_databits_c-1 DOWNTO 0);
          rden_a      : IN STD_LOGIC  := '1';
          rden_b      : IN STD_LOGIC  := '1';
          wren_a      : IN STD_LOGIC  := '0';
          wren_b      : IN STD_LOGIC  := '0';
          q_a         : OUT STD_LOGIC_VECTOR (gpsmem_databits_c-1 DOWNTO 0);
          q_b         : OUT STD_LOGIC_VECTOR (gpsmem_databits_c-1 DOWNTO 0)
        );
      END component gps_ram;

      component ResourceMUX is
        Generic (
          requester_cnt_g       : natural   :=  8 ;
          resource_bits_g       : natural   :=  8 ;
          clock_bitcnt_g        : natural   :=  0 ;
          cross_clock_domain_g  : std_logic := '0'
        ) ;
        Port (
          reset                 : in    std_logic ;
          clk                   : in    std_logic ;
          requesters_in         : in    std_logic_vector (requester_cnt_g-1
                                                              downto 0) ;
          resource_tbl_in       : in    std_logic_2D (requester_cnt_g-1
                                                              downto 0,
                                                      resource_bits_g-1
                                                              downto 0) ;
          receivers_out         : out   std_logic_vector (requester_cnt_g-1
                                                              downto 0) ;
          resources_out         : out   std_logic_vector (resource_bits_g-1
                                                              downto 0)
        ) ;
      end component ResourceMUX ;

      --  GPS Memory access signals.

      signal gpsmem_selected    : std_logic_vector (gpsmem_iobits_c-1
                                                    downto 0) ;

      alias gpsmemdst_addr      : std_logic_vector (gpsmem_addrbits_c-1
                                                    downto 0) is
                                  gpsmem_selected (gpsmem_addrbits_c-1
                                                   downto 0) ;
      alias gpsmemdst_writeto   : std_logic_vector (gpsmem_databits_c-1
                                                    downto 0) is
                                  gpsmem_selected (gpsmem_addrbits_c +
                                                   gpsmem_databits_c - 1
                                                   downto
                                                   gpsmem_addrbits_c) ;
      alias gpsmemdst_read_en   : std_logic is
                                  gpsmem_selected (gpsmem_addrbits_c +
                                                   gpsmem_databits_c) ;
      alias gpsmemdst_write_en  : std_logic is
                                  gpsmem_selected (gpsmem_addrbits_c +
                                                   gpsmem_databits_c + 1) ;
      alias gpsmemdst_clk       : std_logic is
                                  gpsmem_selected (gpsmem_addrbits_c +
                                                   gpsmem_databits_c + 2) ;

    begin

      --  Memory component.  Clock is triggered on negative going edge to
      --  allow input signals to propagate in one half clock cycle and to
      --  produce output by the next clock cycle.  The memory is fast enough
      --  to produce output in less than one half clock cycle.

      gps_ramblocks : gps_ram
        Port Map (
          address_a               => gpsmemsrc_addr,
          address_b               => gpsmemdst_addr,
          clock_a                 => gpsmemsrc_clk,
          clock_b                 => gpsmemdst_clk,
          data_a                  => gpsmemsrc_writeto,
          data_b                  => gpsmemdst_writeto,
          rden_a                  => gpsmemsrc_read_en,
          rden_b                  => gpsmemdst_read_en,
          wren_a                  => gpsmemsrc_write_en,
          wren_b                  => gpsmemdst_write_en,
          q_a                     => gpsmemsrc_readfrom,
          q_b                     => gpsmemdst_readfrom
        ) ;

      --  Resource multiplexer.

      gps_resmux : ResourceMUX
        Generic Map (
          requester_cnt_g         => gpsmemrq_count_c,
          resource_bits_g         => gpsmem_iobits_c,
          clock_bitcnt_g          => 1,
          cross_clock_domain_g    => '1'
        )
        Port Map (
          reset                   => reset,
          clk                     => master_gated_clk,
          requesters_in           => gpsmem_requesters,
          resource_tbl_in         => gpsmem_input_tbl,
          receivers_out           => gpsmem_receivers,
          resources_out           => gpsmem_selected
        ) ;

  end generate use_GPS_RAM ;

  no_use_GPS_RAM:
    if (Collar_Control_useGPSRAM_c = '0') generate

      gpsmemsrc_readfrom        <= (others => '0') ;
      gpsmemdst_readfrom        <= (others => '0') ;
      gpsmem_receivers          <= gpsmem_requesters ;

  end generate no_use_GPS_RAM ;

  --------------------------------------------------------------------------
  --  GPS Message controller.
  --------------------------------------------------------------------------

  use_GPS:
    if (Collar_Control_useGPS_c = '1') generate

      component GPSmessages is

        Generic (
          clk_freq_g            : natural := 50e6 ;
          mem_addrbits_g        : natural := 9 ;
          mem_databits_g        : natural := 8
        ) ;
        Port (
          reset                 : in    std_logic ;
          clk                   : in    std_logic ;
          curtime_in            : in    std_logic_vector (gps_time_bits_c-1
                                                          downto 0) ;
          curtime_latch_in      : in    std_logic ;
          curtime_valid_in      : in    std_logic ;
          curtime_vlatch_in     : in    std_logic ;

          gps_enable_in         : in    std_logic ;
          gps_init_start_in     : in    std_logic ;
          gps_init_done_out     : out   std_logic ;
          pollinterval_in       : in    unsigned (13 downto 0) ;
          datavalid_out         : out   std_logic_vector (msg_ram_blocks_c-1
                                                          downto 0) ;
          gpsmem_clk_out        : out   std_logic ;
          gpsmem_addr_out       : out   std_logic_vector (mem_addrbits_g-1
                                                          downto 0) ;
          gpsmem_read_en_out    : out   std_logic ;
          gpsmem_write_en_out   : out   std_logic ;
          gpsmem_readfrom_in    : in    std_logic_vector (mem_databits_g-1
                                                          downto 0) ;
          gpsmem_writeto_out    : out   std_logic_vector (mem_databits_g-1
                                                          downto 0) ;
          gps_rx_in             : in    std_logic ;
          gps_tx_out            : out   std_logic ;
          timemarker_out        : out   std_logic ;
          gps_timepulse_in      : in    std_logic ;
          aop_running_out       : out   std_logic ;
          busy_out              : out   std_logic
        ) ;
      end component GPSmessages ;

      --  GPS I/O mapping and control signals.

      signal gps_rx           : std_logic ;
      signal gps_tx           : std_logic ;
      signal gps_timemark     : std_logic ;
      signal gps_timepulse    : std_logic ;

      signal poll_int         : unsigned (13 downto 0) :=
                                        TO_UNSIGNED (15, 14) ;

    begin

      gps_ctl : GPSmessages
        Generic Map (
          clk_freq_g            => master_clk_freq_c,
          mem_addrbits_g        => gpsmemsrc_addrbits_c,
          mem_databits_g        => gpsmemsrc_databits_c
        )
        Port Map (
          reset                 => reset,
          clk                   => master_clk,
          curtime_in            => reset_time,
          curtime_latch_in      => systime_latch,
          curtime_valid_in      => systime_valid,
          curtime_vlatch_in     => systime_vlatch,
          gps_enable_in         => CTL_GPS_On,
          gps_init_start_in     => not gps_ready,
          gps_init_done_out     => gps_ready,
          pollinterval_in       => poll_int,
          datavalid_out         => gps_databanks,
          gpsmem_clk_out        => gpsmemsrc_clk,
          gpsmem_addr_out       => gpsmemsrc_addr,
          gpsmem_read_en_out    => gpsmemsrc_read_en,
          gpsmem_write_en_out   => gpsmemsrc_write_en,
          gpsmem_readfrom_in    => gpsmemsrc_readfrom,
          gpsmem_writeto_out    => gpsmemsrc_writeto,
          gps_rx_in             => gps_rx,
          gps_tx_out            => gps_tx,
          timemarker_out        => gps_timemark,
          gps_timepulse_in      => gps_timepulse,
          aop_running_out       => aop_running
        ) ;

      ----------------------------------------------------------------------
      --  All I/O lines forced low when device is off, otherwise they are
      --  driven from the component.
      ----------------------------------------------------------------------

      gps_rx                  <= gps_rx_io ;
      gps_timepulse           <= gps_timepulse_io ;

      gps_on : process (CTL_GPS_On, gps_tx, gps_timemark)
      begin
        if (CTL_GPS_On = '0') then
          gps_rx_io           <= '0' ;
          gps_tx_out          <= '0' ;
          gps_timemark_out    <= '0' ;
          gps_timepulse_io    <= '0' ;
        else
          gps_rx_io           <= 'Z' ;
          gps_tx_out          <= gps_tx ;
          gps_timemark_out    <= gps_timemark ;
          gps_timepulse_io    <= 'Z' ;
        end if ;
      end process gps_on ;

  end generate use_GPS ;

  no_use_GPS:
    if (Collar_Control_useGPS_c = '0') generate

      gps_ready               <= '1' ;

      gps_rx_io               <= '0' ;
      gps_tx_out              <= '0' ;
      gps_timemark_out        <= '0' ;
      gps_timepulse_io        <= '0' ;

      gpsmemsrc_addr          <= (others => '0') ;
      gpsmemsrc_clk           <= '0' ;
      gpsmemsrc_writeto       <= (others => '0') ;
      gpsmemsrc_read_en       <= '0' ;
      gpsmemsrc_write_en      <= '0' ;
      aop_running             <= '0' ;

  end generate no_use_GPS ;

  --------------------------------------------------------------------------
  --  Inertial sensor controller.
  --------------------------------------------------------------------------

  use_Inertial:
    if (Collar_Control_useInertial_c = '1') generate

      component LSM9DS1_top is
        Generic (
          IMU_AXIS_WORD_LENGTH_BYTES  : natural := 2;
          command_used_g              : std_logic := '1';
          address_used_g              : std_logic := '0';
          command_width_bytes_g       : natural := 1;
          address_width_bytes_g       : natural := 1;
          data_length_bit_width_g     : natural := 10
        ) ;
        Port (
          clk                   : in    std_logic ;
          rst_n                 : in    std_logic ;

          startup               : in    std_logic;

          curtime_in            : in    std_logic_vector
                                          (gps_time_bytes_c*8-1 downto 0) ;
          curtime_latch_in      : in    std_logic ;
          curtime_valid_in      : in    std_logic ;
          curtime_vlatch_in     : in    std_logic ;

          gyro_data_rdy   : out     std_logic;
          accel_data_rdy  : out     std_logic;
          mag_data_rdy    : out     std_logic;
          temp_data_rdy   : out     std_logic;

          gyro_data_x     : out     std_logic_vector(IMU_AXIS_WORD_LENGTH_BYTES*8 - 1 downto 0);
          gyro_data_y     : out     std_logic_vector(IMU_AXIS_WORD_LENGTH_BYTES*8 - 1 downto 0);
          gyro_data_z     : out     std_logic_vector(IMU_AXIS_WORD_LENGTH_BYTES*8 - 1 downto 0);

          accel_data_x    : out     std_logic_vector(IMU_AXIS_WORD_LENGTH_BYTES*8 - 1 downto 0);
          accel_data_y    : out     std_logic_vector(IMU_AXIS_WORD_LENGTH_BYTES*8 - 1 downto 0);
          accel_data_z    : out     std_logic_vector(IMU_AXIS_WORD_LENGTH_BYTES*8 - 1 downto 0);

          mag_data_x      : out     std_logic_vector(IMU_AXIS_WORD_LENGTH_BYTES*8 - 1 downto 0);
          mag_data_y      : out     std_logic_vector(IMU_AXIS_WORD_LENGTH_BYTES*8 - 1 downto 0);
          mag_data_z      : out     std_logic_vector(IMU_AXIS_WORD_LENGTH_BYTES*8 - 1 downto 0);

          temp_data       : out     std_logic_vector(IMU_AXIS_WORD_LENGTH_BYTES*8 - 1 downto 0);

          sclk            : out     std_logic;
          mosi            : out     std_logic;
          miso_XL_G       : in      std_logic;
          miso_M          : in      std_logic;
          cs_XL_G         : out     std_logic;
          cs_M            : out     std_logic;

          INT_M           : in      std_logic;
          DRDY_M          : in      std_logic;
          INT1_A_G        : in      std_logic;
          INT2_A_G        : in      std_logic;

          gyro_fpga_time  : out std_logic_vector (gps_time_bytes_c*8-1 downto 0);
          accel_fpga_time : out std_logic_vector (gps_time_bytes_c*8-1 downto 0);
          mag_fpga_time   : out std_logic_vector (gps_time_bytes_c*8-1 downto 0);
          temp_fpga_time  : out std_logic_vector (gps_time_bytes_c*8-1 downto 0)
        ) ;
      end component LSM9DS1_top ;

      --  Inertial module I/O mapping signals.

      signal ms_clock         : std_logic ;
      signal ms_mosi          : std_logic ;
      signal ms_cs_accgyro    : std_logic ;
      signal ms_miso_accgyro  : std_logic ;
      signal ms_int1_accgyro  : std_logic ;
      signal ms_int2_accgyro  : std_logic ;
      signal ms_cs_mag        : std_logic ;
      signal ms_miso_mag      : std_logic ;
      signal ms_int_mag       : std_logic ;
      signal ms_drdy_mag      : std_logic ;

    begin

      im : LSM9DS1_top
        Generic Map (
          IMU_AXIS_WORD_LENGTH_BYTES  => im_datalen_c
        )
        Port Map (
          clk                 => spi_clk,
          rst_n               => (not reset) and CTL_InertialOn1p8 and
                                                 CTL_InertialOn2p5,

          startup             => im_startup,

          curtime_in          => reset_time_bytes,
          curtime_latch_in    => systime_latch,
          curtime_valid_in    => systime_valid,
          curtime_vlatch_in   => systime_vlatch,

          gyro_data_rdy       => im_gyro_data_rdy,
          accel_data_rdy      => im_accel_data_rdy,
          mag_data_rdy        => im_mag_data_rdy,
          temp_data_rdy       => im_temp_data_rdy,

          gyro_data_x         => im_gyro_data_x,
          gyro_data_y         => im_gyro_data_y,
          gyro_data_z         => im_gyro_data_z,

          accel_data_x        => im_accel_data_x,
          accel_data_y        => im_accel_data_y,
          accel_data_z        => im_accel_data_z,

          mag_data_x          => im_mag_data_x,
          mag_data_y          => im_mag_data_y,
          mag_data_z          => im_mag_data_z,

          temp_data           => im_temp_data,

          sclk                => ms_clock,
          mosi                => ms_mosi,
          miso_XL_G           => ms_miso_accgyro,
          miso_M              => ms_miso_mag,
          cs_XL_G             => ms_cs_accgyro,
          cs_M                => ms_cs_mag,

          INT_M               => ms_int_mag,
          DRDY_M              => ms_drdy_mag,
          INT1_A_G            => ms_int1_accgyro,
          INT2_A_G            => ms_int2_accgyro,

          gyro_fpga_time      => im_gyro_time,
          accel_fpga_time     => im_accel_time,
          mag_fpga_time       => im_mag_time,
          temp_fpga_time      => im_temp_time
        ) ;

      ----------------------------------------------------------------------
      --  All I/O lines forced low when device is off, otherwise they are
      --  driven from the component.
      ----------------------------------------------------------------------

      ms_miso_accgyro         <= ms_miso_accgyro_io ;
      ms_int1_accgyro         <= ms_int1_accgyro_io ;
      ms_int2_accgyro         <= ms_int2_accgyro_io ;
      ms_miso_mag             <= ms_miso_mag_io ;
      ms_int_mag              <= ms_int_mag_io ;
      ms_drdy_mag             <= ms_drdy_mag_io ;

      inertial_on : process (CTL_InertialOn1p8, CTL_InertialOn2p5,
                             ms_clock, ms_mosi,
                             ms_cs_accgyro, ms_cs_mag)
      begin
        if (CTL_InertialOn1p8 = '0' or CTL_InertialOn2p5 = '0') then
          ms_clk              <= '0' ;
          ms_mosi_out         <= '0' ;
          ms_cs_accgyro_out   <= '0' ;
          ms_miso_accgyro_io  <= '0' ;
          ms_int1_accgyro_io  <= '0' ;
          ms_int2_accgyro_io  <= '0' ;
          ms_cs_mag_out       <= '0' ;
          ms_miso_mag_io      <= '0' ;
          ms_int_mag_io       <= '0' ;
          ms_drdy_mag_io      <= '0' ;
        else
          ms_clk              <= ms_clock ;
          ms_mosi_out         <= ms_mosi ;
          ms_cs_accgyro_out   <= ms_cs_accgyro ;
          ms_miso_accgyro_io  <= 'Z' ;
          ms_int1_accgyro_io  <= 'Z' ;
          ms_int2_accgyro_io  <= 'Z' ;
          ms_cs_mag_out       <= ms_cs_mag ;
          ms_miso_mag_io      <= 'Z' ;
          ms_int_mag_io       <= 'Z' ;
          ms_drdy_mag_io      <= 'Z' ;
        end if ;
      end process inertial_on ;

    end generate use_Inertial ;

  no_use_Inertial:
    if (Collar_Control_useInertial_c = '0') generate

      ms_clk                  <= '0' ;
      ms_mosi_out             <= '0' ;

      ms_cs_accgyro_out       <= '0' ;
      ms_miso_accgyro_io      <= '0' ;
      ms_int1_accgyro_io      <= '0' ;
      ms_int2_accgyro_io      <= '0' ;

      ms_cs_mag_out           <= '0' ;
      ms_miso_mag_io          <= '0' ;
      ms_int_mag_io           <= '0' ;
      ms_drdy_mag_io          <= '0' ;

      im_gyro_data_rdy        <= '0' ;
      im_accel_data_rdy       <= '0' ;
      im_mag_data_rdy         <= '0' ;
      im_temp_data_rdy        <= '0' ;

      im_gyro_data_x          <= (others => '0') ;
      im_gyro_data_y          <= (others => '0') ;
      im_gyro_data_z          <= (others => '0') ;
      im_accel_data_x         <= (others => '0') ;
      im_accel_data_y         <= (others => '0') ;
      im_accel_data_z         <= (others => '0') ;
      im_mag_data_x           <= (others => '0') ;
      im_mag_data_y           <= (others => '0') ;
      im_mag_data_z           <= (others => '0') ;
      im_temp_data            <= (others => '0') ;

      im_gyro_time            <= (others => '0') ;
      im_accel_time           <= (others => '0') ;
      im_mag_time             <= (others => '0') ;
      im_temp_time            <= (others => '0') ;

    end generate no_use_Inertial ;

  --------------------------------------------------------------------------
  --  Magnetic Memory Buffer
  --------------------------------------------------------------------------

  use_MagMemBuffer:
    if (Collar_Control_useMagMemBuffer_c = '1') generate

      component magmem_ram IS
        PORT
        (
          address_a   : IN STD_LOGIC_VECTOR (magmem_addrbits_c-1 DOWNTO 0);
          address_b   : IN STD_LOGIC_VECTOR (magmem_addrbits_c-1 DOWNTO 0);
          clock_a     : IN STD_LOGIC  := '1';
          clock_b     : IN STD_LOGIC ;
          data_a      : IN STD_LOGIC_VECTOR (magmem_databits_c-1 DOWNTO 0);
          data_b      : IN STD_LOGIC_VECTOR (magmem_databits_c-1 DOWNTO 0);
          rden_a      : IN STD_LOGIC  := '1';
          rden_b      : IN STD_LOGIC  := '1';
          wren_a      : IN STD_LOGIC  := '0';
          wren_b      : IN STD_LOGIC  := '0';
          q_a         : OUT STD_LOGIC_VECTOR (magmem_databits_c-1 DOWNTO 0);
          q_b         : OUT STD_LOGIC_VECTOR (magmem_databits_c-1 DOWNTO 0)
        );
      END component magmem_ram;

      component ResourceMUX is
        Generic (
          requester_cnt_g       : natural   :=  8 ;
          resource_bits_g       : natural   :=  8 ;
          clock_bitcnt_g        : natural   :=  0 ;
          cross_clock_domain_g  : std_logic := '0'
        ) ;
        Port (
          reset                 : in    std_logic ;
          clk                   : in    std_logic ;
          requesters_in         : in    std_logic_vector (requester_cnt_g-1
                                                              downto 0) ;
          resource_tbl_in       : in    std_logic_2D (requester_cnt_g-1
                                                              downto 0,
                                                      resource_bits_g-1
                                                              downto 0) ;
          receivers_out         : out   std_logic_vector (requester_cnt_g-1
                                                              downto 0) ;
          resources_out         : out   std_logic_vector (resource_bits_g-1
                                                              downto 0)
        ) ;
      end component ResourceMUX ;

      --  Magnetic Memory Buffer access signals.

      signal magmem_selected    : std_logic_vector (magmem_iobits_c-1
                                                    downto 0) ;

      alias magmemsrc_addr      : std_logic_vector (magmem_addrbits_c-1
                                                    downto 0) is
                                  magmem_selected (magmem_addrbits_c-1
                                                   downto 0) ;
      alias magmemsrc_writeto   : std_logic_vector (magmem_databits_c-1
                                                    downto 0) is
                                  magmem_selected (magmem_addrbits_c +
                                                   magmem_databits_c - 1
                                                   downto
                                                   magmem_addrbits_c) ;
      alias magmemsrc_read_en   : std_logic is
                                  magmem_selected (magmem_addrbits_c +
                                                   magmem_databits_c) ;
      alias magmemsrc_write_en  : std_logic is
                                  magmem_selected (magmem_addrbits_c +
                                                   magmem_databits_c + 1) ;
      alias magmemsrc_clk       : std_logic is
                                  magmem_selected (magmem_addrbits_c +
                                                   magmem_databits_c + 2) ;

    begin

      magmem_buff_busy  <= '1' when ((unsigned (magmem_requesters) /= 0)  or
                                     (unsigned (magmem_receivers)  /= 0))
                               else '0' ;

      --  Memory component.  Clock is triggered on negative going edge to
      --  allow input signals to propagate in one half clock cycle and to
      --  produce output by the next clock cycle.  The memory is fast enough
      --  to produce output in less than one half clock cycle.

      magmem_ramblocks : magmem_ram
        Port Map (
          address_a               => magmemsrc_addr,
          address_b               => magmemdst_addr,
          clock_a                 => magmemsrc_clk,
          clock_b                 => magmemdst_clk,
          data_a                  => magmemsrc_writeto,
          data_b                  => magmemdst_writeto,
          rden_a                  => magmemsrc_read_en,
          rden_b                  => magmemdst_read_en,
          wren_a                  => magmemsrc_write_en,
          wren_b                  => magmemdst_write_en,
          q_a                     => magmemsrc_readfrom,
          q_b                     => magmemdst_readfrom
        ) ;

      --  Resource multiplexer.

      magmem_resmux : ResourceMUX
        Generic Map (
          requester_cnt_g         => magmemrq_count_c,
          resource_bits_g         => magmem_iobits_c,
          clock_bitcnt_g          => 1,
          cross_clock_domain_g    => '1'
        )
        Port Map (
          reset                   => reset,
          clk                     => master_gated_clk,
          requesters_in           => magmem_requesters,
          resource_tbl_in         => magmem_input_tbl,
          receivers_out           => magmem_receivers,
          resources_out           => magmem_selected
        ) ;

  end generate use_MagMemBuffer ;

  no_use_MagMemBuffer:
    if (Collar_Control_useMagMemBuffer_c = '0') generate

      magmemsrc_readfrom        <= (others => '0') ;
      magmemdst_readfrom        <= (others => '0') ;
      magmem_receivers          <= magmem_requesters ;

      magmem_buff_busy          <= '0' ;

  end generate no_use_MagMemBuffer ;

  --------------------------------------------------------------------------
  --  Magnetic RAM control.
  --------------------------------------------------------------------------

  use_Magmem:
    if (Collar_Control_useMagMem_c = '1') generate

      component magmem_controller is
        Generic (
          clk_freq_g              : natural := 50E6;
          mag_interval_ms_g       : natural := 2;
          tRDP_sleep_mode_exit_time_us  : natural := 2;
          buffer_bytes_g          : natural := 1024;
          buffer_num_g            : natural := 2;

          command_used_g          : std_logic := '1';
          address_used_g          : std_logic := '1';
          command_width_bytes_g   : natural := 1;
          address_width_bytes_g   : natural := 3;
          data_length_bit_width_g : natural := 10
        ) ;
        Port (
          clk               : in  std_logic ;
          rst_n             : in  std_logic ;

          startup           : in  std_logic;
          startup_finished  : out std_logic;
          mag_ram_clk_a     : out std_logic;
          mag_ram_wr_en_a   : out std_logic;
          mag_ram_rd_en_a   : out std_logic;
          mag_ram_address_a : out std_logic_vector(natural(trunc(log2(real(buffer_bytes_g-1)))) downto 0);
          mag_ram_data_a    : out std_logic_vector(7 downto 0);

          mem_req_a_out     : out std_logic;
          mem_rec_a_in      : in std_logic;

          ram_mag_q_b       : in std_logic_vector(7 downto 0);
          ram_mag_data_b    : out std_logic_vector(7 downto 0);
          mag_ram_clk_b     : out std_logic;
          mag_ram_rd_en_b   : out std_logic;
          mag_ram_wr_en_b   : out std_logic;
          mag_ram_address_b : out std_logic_vector(natural(trunc(log2(real(buffer_bytes_g-1)))) downto 0);

          miso              : in std_logic;
          mosi              : out std_logic;
          sclk              : out std_logic;
          cs_n              : out std_logic;

          fpga_time         : in  std_logic_vector(gps_time_bits_c-1 downto 0);
          current_active_ram_buffer : out   std_logic_vector(natural(trunc(log2(real(
                                        buffer_num_g-1)))) downto 0)
        ) ;
      end component magmem_controller ;

      --  Magnetic Memory I/O mapping signals.

      signal magmem_clock       : std_logic ;
      signal magmem_cs          : std_logic ;
      signal magmem_mosi        : std_logic ;
      signal magmem_miso        : std_logic ;

      --  Magnetic Memory source access signals.

      signal magmemsrc_clk      : std_logic ;
      signal magmemsrc_write_en : std_logic ;
      signal magmemsrc_read_en  : std_logic ;
      signal magmemsrc_addr     : std_logic_vector (magmem_addrbits_c-1
                                                    downto 0) ;
      signal magmemsrc_writeto  : std_logic_vector (magmem_databits_c-1
                                                    downto 0) ;
      signal magmemsrc_control  : std_logic_vector (magmem_iobits_c-1
                                                    downto 0) ;

    begin

      magmem : magmem_controller
        Generic Map (
          clk_freq_g        => spi_clk_freq_c,
          buffer_bytes_g    => mm_buffbytes_c,
          buffer_num_g      => mm_buffnum_c
        )
        Port Map (
          clk               => spi_clk,
          rst_n             => (not reset) and CTL_MagMemOn,
          startup           => mm_startup,
          startup_finished  => mm_startup_done,
          mag_ram_clk_a     => magmemsrc_clk,
          mag_ram_wr_en_a   => magmemsrc_write_en,
          mag_ram_rd_en_a   => magmemsrc_read_en,
          mag_ram_address_a => magmemsrc_addr,
          mag_ram_data_a    => magmemsrc_writeto,
          mem_req_a_out     => magmem_requesters (magmemrq_magmem_c),
          mem_rec_a_in      => magmem_receivers  (magmemrq_magmem_c),
          ram_mag_q_b       => magmemdst_readfrom,
          ram_mag_data_b    => magmemdst_writeto,
          mag_ram_clk_b     => magmemdst_clk,
          mag_ram_rd_en_b   => magmemdst_read_en,
          mag_ram_wr_en_b   => magmemdst_write_en,
          mag_ram_address_b => magmemdst_addr,
          miso              => magmem_miso,
          mosi              => magmem_mosi,
          sclk              => magmem_clock,
          cs_n              => magmem_cs,
          fpga_time         => reset_time,
          current_active_ram_buffer   => mm_buffno
        ) ;

      magmemsrc_control     <= spi_gated_inv_clk  &
                               magmemsrc_write_en & magmemsrc_read_en &
                               magmemsrc_writeto  & magmemsrc_addr ;

      set2D_element (magmemrq_magmem_c, magmemsrc_control,
                     magmem_input_tbl) ;

      ----------------------------------------------------------------------
      --  All I/O lines forced low when device is off, otherwise they are
      --  driven from the component.
      ----------------------------------------------------------------------

      magmem_miso               <= magram_miso_io ;
      magram_writeprot_out      <= '0' ;

      magmem_on : process (CTL_MagMemOn, magmem_clock, magmem_cs,
                           magmem_mosi)
      begin
        if (CTL_MagMemOn = '0') then
          magram_clk            <= '0' ;
          magram_cs_out         <= '0' ;
          magram_mosi_out       <= '0' ;
          magram_miso_io        <= '0' ;
        else
          magram_clk            <= magmem_clock ;
          magram_cs_out         <= magmem_cs ;
          magram_mosi_out       <= magmem_mosi ;
          magram_miso_io        <= 'Z' ;
        end if ;
      end process magmem_on ;

    end generate use_Magmem ;

  no_use_MagMem:
    if (Collar_Control_useMagMem_c = '0') generate

      mm_startup_done         <= '1' ;

      magram_clk              <= '0' ;
      magram_cs_out           <= '0' ;
      magram_mosi_out         <= '0' ;
      magram_miso_io          <= '0' ;
      magram_writeprot_out    <= '0' ;

      magmemdst_writeto       <= (others => '0') ;
      magmemdst_read_en       <= '0' ;
      magmemdst_write_en      <= '0' ;
      magmemdst_addr          <= (others => '0') ;

      magmem_requesters (magmemrq_magmem_c)  <= '0' ;

      end generate no_use_MagMem ;

  --------------------------------------------------------------------------
  --  Microphone control.
  --------------------------------------------------------------------------

  use_PDMmic:
    if (Collar_Control_usePDMmic_c = '1') generate

      component mems_top_16 is
        port (
          clk         :   IN    std_logic;
          rst_n       :   IN    std_logic;
          clk_enable  :   IN    std_logic;
          pdm_bit     :   IN    std_logic;
          filter_out  :   OUT   std_logic_vector(15 DOWNTO 0); -- sfix16
          clock_out   :   OUT   std_logic  --clk / 64.
          );
      end component mems_top_16;

      --  Microphone I/O mapping signals.

      signal mic_clock    : std_logic ;
      signal mic_right    : std_logic ;
      signal mic_left     : std_logic ;

      -- Microphone Test Signals
      signal mic_left_sample_clk_f  : std_logic;

    begin

      --  The microphones will use the SPI clock as their driver.

      mic_clock           <= spi_clk ;

      mright : mems_top_16
        port map (
          clk             => mic_clock,
          rst_n           => (not reset) and CTL_MicRightOn,
          clk_enable      => '1',
          pdm_bit         => mic_right,
          filter_out      => mic_right_sample,
          clock_out       => mic_right_sample_clk
        ) ;

      mleft : mems_top_16
        port map (
          clk             => mic_clock,
          rst_n           => (not reset) and CTL_MicLeftOn,
          clk_enable      => '1',
          pdm_bit         => mic_left,
          --filter_out      => mic_left_sample,
          clock_out       => mic_left_sample_clk
        ) ;

      ----------------------------------------------------------------------
      --  All I/O lines forced low when device is off, otherwise they are
      --  driven from the component.
      ----------------------------------------------------------------------

      mic_right                 <= mic_right_io ;
      mic_left                  <= mic_left_io ;

      mics_on : process (CTL_MicLeftOn, CTL_MicRightOn, mic_clock)
      begin
        if (CTL_MicLeftOn = '0' and CTL_MicRightOn = '0') then
          mic_clk               <= '0' ;
          mic_left_io           <= '0' ;
          mic_right_io          <= '0' ;
        else
          mic_clk               <= mic_clock ;

          if (CTL_MicLeftOn = '0') then
            mic_left_io         <= '0' ;
          else
            mic_left_io         <= 'Z' ;
          end if ;

          if (CTL_MicRightOn = '0') then
            mic_right_io        <= '0' ;
          else
            mic_right_io        <= 'Z' ;
          end if ;
        end if ;
      end process mics_on ;



      --TEST PROCESS
      mems_mic_counter:  process(mic_clock, reset)
      begin
      if (reset = '1') then
        mic_left_sample   <= (others => '0');
        mic_left_sample_clk_f <= '0';
      elsif (mic_clock'event and mic_clock = '1') then
        if (mic_left_sample_clk_f /= mic_left_sample_clk ) then
          mic_left_sample_clk_f <= mic_left_sample_clk;
          if (mic_left_sample_clk = '1') then
            mic_left_sample <= std_logic_vector(unsigned(mic_left_sample) + 1);
          end if;
        end if;
      end if;
      end process;
      --TEST PROCESS

    end generate use_PDMmic ;

  no_use_PDMmic:
    if (Collar_Control_usePDMmic_c = '0') generate

      mic_clk                 <= '0' ;
      mic_left_io             <= '0' ;
      mic_right_io            <= '0' ;

      mic_left_sample         <= (others => '0') ;
      mic_left_sample_clk     <= '0' ;

      mic_right_sample        <= (others => '0') ;
      mic_right_sample_clk    <= '0' ;

    end generate no_use_PDMmic ;

  --------------------------------------------------------------------------
  --  Radio control.
  --------------------------------------------------------------------------

  use_Radio:
    if (Collar_Control_useRadio_c = '1') generate

      --  Radio I/O mapping signals.

      signal radio_clock      : std_logic ;
      signal radio_data       : std_logic_vector (radio_data_io'length-1
                                                  downto 0) ;

    begin

      --  The radio will run at SPI speed.

      radio_clock               <= spi_clk ;

      ----------------------------------------------------------------------
      --  All I/O lines forced low when device is off, otherwise they are
      --  driven from the component.
      ----------------------------------------------------------------------

      radio_data                <= radio_data_io ;

      radio_on : process (CTL_DataTX_On, radio_clock)
      begin
        if (CTL_DataTX_On = '0') then
          radio_clk             <= '0' ;
          radio_data_io         <= (others => '0') ;
        else
          radio_clk             <= radio_clock ;
          radio_data_io         <= (others => 'Z') ;
        end if ;
      end process radio_on ;

    end generate use_Radio ;

  no_use_Radio:
    if (Collar_Control_useRadio_c = '0') generate

      radio_clk               <= '0' ;
      radio_data_io           <= (others => '0') ;

    end generate no_use_Radio ;

  --------------------------------------------------------------------------
  --  Flash Block
  --------------------------------------------------------------------------

  use_FlashBlock:
    if (Collar_Control_useFlashBlock_c = '1') generate

      component FlashBlock is

        Generic (
          fpga_time_length_bytes_g  : natural := 9;
          time_bytes_g              : natural := 9 ;
          event_bytes_g             : natural := 2 ;

          rtc_time_bytes_g          : natural := 4;
          num_mics_active_g         : natural := 1;

          counter_data_size_g       : natural     := 8 ;
          counter_address_size_g    : natural     := 9 ;
          counters_g                : natural     := 10 ;

          gps_buffer_bytes_g            : natural := 512;
          imu_axis_word_length_bytes_g  : natural := 2;
          sdram_input_buffer_bytes_g    : natural := 4096;
          audio_word_bytes_g            : natural := 2
      ) ;
        Port (
          clock_sys             : in    std_logic ;
          rst_n                 : in    std_logic ;
          clk_enable            : in    std_logic;

          log_status            : in    std_logic ;

          curtime_in            : in    std_logic_vector
                                          (gps_time_bytes_c*8-1 downto 0) ;
          curtime_latch_in      : in    std_logic ;
          curtime_valid_in      : in    std_logic ;
          curtime_vlatch_in     : in    std_logic ;
          log_events            : in    std_logic;

          gyro_data_rdy   : in    std_logic;
          accel_data_rdy  : in    std_logic;
          mag_data_rdy    : in    std_logic;
          temp_data_rdy   : in    std_logic;


          gyro_data_x     :in     std_logic_vector(
                                  imu_axis_word_length_bytes_g*8 - 1 downto 0);
          gyro_data_y     :in     std_logic_vector(
                                  imu_axis_word_length_bytes_g*8 - 1 downto 0);
          gyro_data_z     :in     std_logic_vector(
                                  imu_axis_word_length_bytes_g*8 - 1 downto 0);

          accel_data_x    :in     std_logic_vector(
                                  imu_axis_word_length_bytes_g*8 - 1 downto 0);
          accel_data_y    :in     std_logic_vector(
                                  imu_axis_word_length_bytes_g*8 - 1 downto 0);
          accel_data_z    :in     std_logic_vector(
                                  imu_axis_word_length_bytes_g*8 - 1 downto 0);

          mag_data_x      :in     std_logic_vector(
                                  imu_axis_word_length_bytes_g*8 - 1 downto 0);
          mag_data_y      :in     std_logic_vector(
                                  imu_axis_word_length_bytes_g*8 - 1 downto 0);
          mag_data_z      :in     std_logic_vector(
                                  imu_axis_word_length_bytes_g*8 - 1 downto 0);

          temp_data       :in     std_logic_vector(
                                  imu_axis_word_length_bytes_g*8 - 1 downto 0);

          audio_data_rdy          : in std_logic;
          audio_data              : in std_logic_vector(
                                    audio_word_bytes_g*8  - 1 downto 0);

          flashblock_inbuf_data       : out    std_logic_vector(7 downto 0);
          flashblock_inbuf_wr_en      : out    std_logic;
          flashblock_inbuf_clk        : out    std_logic;
          flashblock_inbuf_addr       : out   std_logic_vector(
                                              natural(trunc(log2(real(
                                              sdram_input_buffer_bytes_g-1))))
                                              downto 0);

          flashblock_gpsbuf_addr      : out   std_logic_vector(
                                              natural(trunc(log2(real(
                                              gps_buffer_bytes_g-1))))
                                              downto 0);
          flashblock_gpsbuf_rd_en     : out   std_logic;
          flashblock_gpsbuf_clk       : out   std_logic;
          gpsbuf_flashblock_data      : in    std_logic_vector(7 downto 0);

          gps_req_out       : out   std_logic;
          gps_rec_in        : in    std_logic;


          posbank     :in std_logic;
          tmbank      :in std_logic;

          gyro_fpga_time  :in std_logic_vector (gps_time_bytes_c*8-1 downto 0);
          accel_fpga_time :in std_logic_vector (gps_time_bytes_c*8-1 downto 0);
          mag_fpga_time :in std_logic_vector (gps_time_bytes_c*8-1 downto 0);
          temp_fpga_time :in std_logic_vector (gps_time_bytes_c*8-1 downto 0);

          rtc_time_in : in std_logic_vector (rtc_time_bytes_g*8-1 downto 0);

          flashblock_counter_rd_wr_addr  : out   std_logic_vector(
                                              counter_address_size_g-1 downto 0);
          flashblock_counter_rd_en    : out   std_logic;
          flashblock_counter_wr_en    : out   std_logic;
          flashblock_counter_clk      : out   std_logic;
          flashblock_counter_lock     : out   std_logic;
          flashblock_counter_data     : out   std_logic_vector(
                                              counter_data_size_g-1 downto 0);
          counter_flashblock_data     : in    std_logic_vector(
                                              counter_data_size_g-1 downto 0);

          flashblock_sdram_2k_accumulated : out  std_logic;

          mem_req_a_out           : out std_logic;
          mem_rec_a_in            : in std_logic;

          fb_magram_clk_a_out     : out std_logic;
          fb_magram_wr_en_a_out   : out std_logic;
          fb_magram_rd_en_a_out   : out std_logic;
          fb_magram_address_a_out : out std_logic_vector(natural(trunc(log2(real(
                                      (magmem_buffer_bytes/magmem_buffer_num)-1)))) downto 0);
          fb_magram_data_a_out    : out std_logic_vector(7 downto 0);
          magram_fb_q_a_in        : in std_logic_vector(7 downto 0);


          force_wr_en             : out  std_logic;
          sdram_empty_in          : in   std_logic;

          crit_event              : in   std_logic;
          blocks_past_crit        : out  std_logic_vector(7 downto 0)
      ) ;

      end component FlashBlock ;


      --  Flash Block to GPS Memory communications signals.

      signal fb_gpsmem_clk        : std_logic ;
      signal fb_gpsmem_rd_en      : std_logic ;
      signal fb_gpsmem_addr       : std_logic_vector (gpsmem_addrbits_c-1
                                                      downto 0) ;
      signal fb_gpsmem_control    : std_logic_vector (gpsmem_iobits_c-1
                                                      downto 0) ;

      --  Flash Block to Magnetic Memory communications signals.

      signal fb_magmem_clk        : std_logic ;
      signal fb_magmem_wr_en      : std_logic ;
      signal fb_magmem_rd_en      : std_logic ;
      signal fb_magmem_addr       : std_logic_vector(natural(trunc(log2(
                                    real((magmem_buffer_bytes/magmem_buffer_num)-1)
                                    ))) downto 0);
      -- signal fb_magmem_addr       : std_logic_vector (magmem_addrbits_c-1
                                                      -- downto 0) ;
      signal fb_magmem_writeto    : std_logic_vector (magmem_databits_c-1
                                                      downto 0) ;
      signal fb_magmem_control    : std_logic_vector (magmem_iobits_c-1
                                                      downto 0) ;

      --  The audio data from the microphones is concatinated into a single
      --  word.

      constant audio_bytes_c  : natural :=
          natural (trunc (real (mic_left_sample'length +
                                mic_right_sample'length - 1) / 8.0)) + 1 ;

      signal audio_word       : std_logic_vector (audio_bytes_c*8-1
                                                  downto 0) :=
                                                      (others => '0') ;

    begin

      audio_word (mic_left_sample'length +
                  mic_right_sample'length - 1
                  downto 0)                     <= mic_left_sample &
                                                   mic_right_sample ;

      flashblk : FlashBlock
        Generic Map (
          fpga_time_length_bytes_g      => gps_time_bytes_c,
          time_bytes_g                  => gps_time_bytes_c,
          event_bytes_g                 => eventcnt_bytes_c,
          rtc_time_bytes_g              => rtc_time_bytes_c,
          num_mics_active_g             => 2,
          counter_data_size_g         => eventcnt_databits_c,
          counter_address_size_g      => eventcnt_addrbits_c,
          counters_g                  => eventcnt_events_c,
          gps_buffer_bytes_g            => gpsmem_bytecnt_c,
          imu_axis_word_length_bytes_g  => im_datalen_c,
          sdram_input_buffer_bytes_g    => inmem_bytecnt_c,
          audio_word_bytes_g            => 2
        )
        Port Map (
          clock_sys                   => spi_clk,
          rst_n                       => (not reset),
          clk_enable                  => '1',
          log_status                  => SDLogging_status,
          curtime_in                  => reset_time_bytes,
          curtime_latch_in            => systime_latch,
          curtime_valid_in            => systime_valid,
          curtime_vlatch_in           => systime_vlatch,
          log_events                  => eventcnt_changed,
          gyro_data_rdy               => im_gyro_data_rdy,
          accel_data_rdy              => im_accel_data_rdy,
          mag_data_rdy                => im_mag_data_rdy,
          temp_data_rdy               => im_temp_data_rdy,
          gyro_data_x                 => im_gyro_data_x,
          gyro_data_y                 => im_gyro_data_y,
          gyro_data_z                 => im_gyro_data_z,
          accel_data_x                => im_accel_data_x,
          accel_data_y                => im_accel_data_y,
          accel_data_z                => im_accel_data_z,
          mag_data_x                  => im_mag_data_x,
          mag_data_y                  => im_mag_data_y,
          mag_data_z                  => im_mag_data_z,
          temp_data                   => im_temp_data,
          audio_data_rdy              => mic_left_sample_clk,
          audio_data                  => mic_left_sample,
          flashblock_inbuf_data       => sdram_inwr_data,
          flashblock_inbuf_wr_en      => sdram_inwr_en,
          flashblock_inbuf_clk        => sdram_inwr_clk,
          flashblock_inbuf_addr       => sdram_inwr_addr,
          flashblock_gpsbuf_addr      => fb_gpsmem_addr,
          flashblock_gpsbuf_rd_en     => fb_gpsmem_rd_en,
          flashblock_gpsbuf_clk       => fb_gpsmem_clk,
          gpsbuf_flashblock_data      => gpsmemdst_readfrom,
          gps_req_out                 => gpsmem_requesters (gpsmemrq_flashblk_c),
          gps_rec_in                  => gpsmem_receivers (gpsmemrq_flashblk_c),
          posbank                     =>
                            gps_databanks (msg_ubx_nav_sol_ramblock_c),
          tmbank                      =>
                            gps_databanks (msg_ubx_tim_tm2_ramblock_c),
          gyro_fpga_time              => im_gyro_time,
          accel_fpga_time             => im_accel_time,
          mag_fpga_time               => im_mag_time,
          temp_fpga_time              => im_temp_time,
          rtc_time_in                 =>
                            std_logic_vector (rtc_running_seconds),
          flashblock_counter_rd_wr_addr  => evmemdst_addr,
          flashblock_counter_rd_en    => evmemdst_read_en,
          flashblock_counter_wr_en    => evmemdst_write_en,
          flashblock_counter_clk      => evmemdst_clk,
          flashblock_counter_lock     => eventcnt_lock,
          flashblock_counter_data     => evmemdst_writeto,
          counter_flashblock_data     => evmemdst_readfrom,
          flashblock_sdram_2k_accumulated   => sdram_inready,
          mem_req_a_out              =>
                    magmem_requesters (magmemrq_flashblk_c),
          mem_rec_a_in               =>
                  magmem_receivers  (magmemrq_flashblk_c),
          fb_magram_clk_a_out         =>  fb_magmem_clk,
          fb_magram_wr_en_a_out            => fb_magmem_wr_en,
          fb_magram_rd_en_a_out            => fb_magmem_rd_en,
          fb_magram_address_a_out          => fb_magmem_addr,
          fb_magram_data_a_out             => fb_magmem_writeto,
          magram_fb_q_a_in              => magmemsrc_readfrom,

          force_wr_en                 => sdram_forceout,
          sdram_empty_in              => sdram_empty,
          crit_event                  => SDLogging_flush,
          blocks_past_crit            => sdcard_critpast
        ) ;

      fb_gpsmem_control    <= spi_gated_inv_clk   &
                              gpsmem_wren_none_c  & fb_gpsmem_rd_en &
                              gpsmem_wrto_none_c  & fb_gpsmem_addr ;

      set2D_element (gpsmemrq_flashblk_c, fb_gpsmem_control,
                     gpsmem_input_tbl) ;

      fb_magmem_control    <= spi_gated_inv_clk &
                              fb_magmem_wr_en   & fb_magmem_rd_en &
                              fb_magmem_writeto & mm_buffno &
                              fb_magmem_addr ;

      set2D_element (magmemrq_flashblk_c, fb_magmem_control,
                     magmem_input_tbl) ;

    end generate use_FlashBlock ;

  no_use_FlashBlock:
    if (Collar_Control_useFlashBlock_c = '0') generate
      signal fb_gpsmem_control      : std_logic_vector (gpsmem_iobits_c-1
                                                          downto 0) :=
                                            (others => '0') ;
      signal fb_magmem_control      : std_logic_vector (magmem_iobits_c-1
                                                          downto 0) :=
                                            (others => '0') ;
    begin
      gpsmem_requesters (gpsmemrq_flashblk_c) <= '0' ;

      fb_gpsmem_control (gpsmem_iobits_c-1)   <= spi_gated_inv_clk ;
      set2D_element (gpsmemrq_flashblk_c, fb_gpsmem_control,
                     gpsmem_input_tbl) ;

      magmem_requesters (magmemrq_flashblk_c) <= '0' ;

      fb_magmem_control (magmem_iobits_c-1)   <= spi_gated_inv_clk ;
      set2D_element (magmemrq_flashblk_c, fb_magmem_control,
                     magmem_input_tbl) ;

    end generate no_use_FlashBlock ;

  --------------------------------------------------------------------------
  --  Reset occurs on power up or button press of the reset button.
  --------------------------------------------------------------------------

  global_reset : GlobalClock
    Port Map
    (
      ena       => '1',
      inclk     => (not power_up) or reset_pushed,
      outclk    => reset
    ) ;

  reset_poweron : process (master_clk)
  begin
    if (rising_edge (master_clk)) then
      if (pu_counter = pu_count_c) then
        power_up            <= '1' ;
      else
        pu_counter          <= pu_counter + 1 ;
      end if ;
    end if ;
  end process reset_poweron ;

  --  Debounce the reset button by making sure it is held up or down for a
  --  long period of time.

  reset_pb : process (master_clk)
  begin
    if (rising_edge (master_clk)) then

      if (buttons_in (reset_button_c) /= reset_pushed) then
        if (pb_counter = pb_count_c) then
          reset_pushed      <= buttons_in (reset_button_c) ;
          pb_counter        <= (others => '0') ;
        else
          pb_counter        <= pb_counter + 1 ;
        end if ;
      else
        pb_counter          <= (others => '0') ;
      end if ;
    end if ;
  end process reset_pb ;


end architecture structural ;
