----------------------------------------------------------------------------
--
--! @file       PowerController.vhd
--! @brief      Power Controller Top Level.
--! @details    Instanciates and connects all the components that make up
--!             the Power Controller CPLD implementation.
--! @author     Emery Newlon
--! @date       September 2014
--! @copyright  Copyright (C) 2014 Ross K. Snider and Emery L. Newlon
--
--  This program is free software: you can redistribute it and/or modify
--  it under the terms of the GNU General Public License as published by
--  the Free Software Foundation, either version 3 of the License, or
--  (at your option) any later version.
--
--  This program is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--  GNU General Public License for more details.
--
--  You should have received a copy of the GNU General Public License
--  along with this program.  If not, see <http://www.gnu.org/licenses/>.
--
--  Emery Newlon
--  Electrical and Computer Engineering
--  Montana State University
--  610 Cobleigh Hall
--  Bozeman, MT 59717
--  emery.newlon@msu.montana.edu
--
----------------------------------------------------------------------------

library IEEE ;                      --! Use standard library.
use IEEE.STD_LOGIC_1164.ALL ;       --! Use standard logic elements.
use IEEE.NUMERIC_STD.ALL ;          --! Use numeric standard.
use IEEE.MATH_REAL.ALL ;            --! Real number functions.

library GENERAL ;                   --! General libraries
use GENERAL.UTILITIES_PKG.ALL ;

library WORK ;                      --! Local Libaries
use WORK.PC_STATUSCONTROL_PKG.All ;


----------------------------------------------------------------------------
--
--! @brief      Power Controller Top Level.
--! @details    Instanciates and connects all the components that make up
--!             the Power Controller CPLD implementation.
--!
--! @param      master_clk_freq_g Frequency of the system clock in cycles
--!                               per second.
--! @param      master_clk        Clock generated by the system that drives
--!                               everything else.
--! @param      master_clk_out    Output of the master clock to the FPGA.
--!
--! @param      flash_clk_out         Flash clock.
--! @param      flash_cs_out          Flash chip select.
--! @param      pfl_flash_data_io     Parallel Flash Loader Flash data bus.
--! @param      fpga_flash_data_io    FPGA Flash data bus.
--! @param      fpga_toflash_clk_in   FPGA to Flash clock.
--! @param      fpga_toflash_cs_in    FPGA to Flash chip select.
--! @param      fpga_toflash_data_io  FPGA to Flash data bus.
--! @param      fpga_toflash_dir_in   FPGA to Flash data direction.
--!
--! @param      fpga_cnf_dclk_out     FPGA Configuration data clock.
--! @param      fpga_cnf_data_out     FPGA Configuration data to FPGA.  Must
--!                                   not be left floating after
--!                                   configuration.
--! @param      fpga_cnf_nstatus_in   FPGA Configuration status not.  Must
--!                                   have a pull-up resistor.
--! @param      fpga_cnf_conf_done_in FPGA Configuration config done.  Must
--!                                   have a pull-up resistor.
--! @param      fpga_cnf_init_done_in FPGA Configuration init done.  Must
--!                                   have a pull-up resistor.
--! @param      fpga_cnf_nconfig_out  FPGA Configuration configure not.
--!                                   Must have a pull-up resistor if used
--!                                   as an open drain pin.
--!
--! @param      statchg_out       The status register has changed.
--! @param      spi_clk_in        The PC status register / FPGA control
--!                               register SPI bus clock.
--! @param      spi_cs_in         The PC SPI bus chip select.  An SPI
--!                               transfer is initiated when it goes low.
--! @param      spi_mosi_in       Master Out/Slave In SPI data line.
--! @param      spi_miso_out      Master In/Slave Out SPI data line.
--!
--! @param      i2c_clk_io        I2C bus clock is input or output depending
--!                               on the device driving it.
--! @param      i2c_data_io       I2C bus data is driven by the same device
--!                               that is driving the clock.
--!
--! @param      bat_power_out     Battery power switch.
--! @param      bat_recharge_out  Battery recharge switch.
--! @param      bat_int_in        Battery monitor interrupt.
--! @param      bat_int_fpga_out  Battery monitor interrupt to FPGA.
--! @param      bat_low_in        Battery monitor battery low.
--! @param      bat_good_in       Battery monitor battery good.
--!
--! @param      pwr_1p1_run_out   Power on the 1.1 V power supply.
--! @param      pwr_1p1_good_in   The 1.1 V power supply is operating.
--! @param      pwr_2p5_run_out   Power on the 2.5 V power supply.
--! @param      pwr_2p5_good_in   The 2.5 V power supply is operating.
--! @param      pwr_3p3_run_out   Power on the 3.3 V power supply.
--! @param      pwr_3p3_good_in   The 3.3 V power supply is operating.
--! @param      pwr_pwm_out       Use PWM or burst mode.
--!
--! @param      pwr_drive_out     Drive the power switch buffer signals.
--! @param      pwr_clock_out     Power on the clock.
--! @param      pwr_fpga_out      Power on the FPGA 1.8, 2.5, & 3.3 Vcc.
--! @param      pwr_sdram_out     Power on the SDRAM.
--! @param      pwr_mram_out      Power on the Magnetic RAM.
--! @param      pwr_im_out        Power on the Inertial Modules.
--! @param      pwr_gps_out       Power on the GPS.
--! @param      pwr_datatx_out    Power on the Data Transmitter.
--! @param      pwr_micR_out      Power on the Right Hand Microphone.
--! @param      pwr_micL_out      Power on the Left Hand Microphone.
--! @param      pwr_sdcard_out    Power on the SD Cards.
--! @param      pwr_ls_1p8_out    Power on the 1.8 V Level Shifter.
--! @param      pwr_ls_3p3_out    Power on the 3.3 V Level Shifter.
--!
--! @param      solar_max_in      Solar Controller voltage level is at max.
--! @param      solar_on_in       Solar Controller is operating.
--! @param      solar_run_out     Solar Controller is turned on.
--!
--! @param      forced_start_in   A forced startup has been initiated.
--! @param      fpga_fs_out       Forced startup passed to the FPGA.
--! @param      rtc_alarm_in      Alarm interrupt from the Real Time Clock.
--
----------------------------------------------------------------------------

entity PowerController is

  Generic (
    master_clk_freq_g     : natural   := 10e6
  ) ;
  Port (
    master_clk            : in    std_logic ;
    master_clk_out        : out   std_logic ;

    flash_clk_out         : out   std_logic ;
    flash_cs_out          : out   std_logic ;
    pfl_flash_data_io     : inout std_logic_vector (3 downto 0) ;
    fpga_flash_data_io    : inout std_logic_vector (3 downto 0) ;
    fpga_toflash_clk_in   : inout std_logic ;
    fpga_toflash_cs_in    : inout std_logic ;
    fpga_toflash_data_io  : inout std_logic_vector (3 downto 0) ;
    fpga_toflash_dir_in   : inout std_logic ;

    fpga_cnf_dclk_out     : out   std_logic ;
    fpga_cnf_data_out     : out   std_logic ;
    fpga_cnf_nstatus_in   : in    std_logic ;
    fpga_cnf_conf_done_in : in    std_logic ;
    fpga_cnf_init_done_in : in    std_logic ;
    fpga_cnf_nconfig_out  : out   std_logic ;

    statchg_out           : out   std_logic ;
    spi_clk_in            : inout std_logic ;
    spi_cs_in             : inout std_logic ;
    spi_mosi_in           : inout std_logic ;
    spi_miso_out          : out   std_logic ;

    i2c_clk_io            : inout std_logic ;
    i2c_data_io           : inout std_logic ;

    bat_power_out         : out   std_logic ;
    bat_recharge_out      : out   std_logic ;
    bat_int_in            : in    std_logic ;
    bat_int_fpga_out      : inout std_logic ;
    bat_low_in            : in    std_logic ;
    bat_good_in           : in    std_logic ;

    pwr_1p1_run_out       : out   std_logic ;
    pwr_1p1_good_in       : in    std_logic ;
    pwr_2p5_run_out       : out   std_logic ;
    pwr_2p5_good_in       : in    std_logic ;
    pwr_3p3_run_out       : out   std_logic ;
    pwr_3p3_good_in       : in    std_logic ;
    pwr_pwm_out           : out   std_logic ;

    pwr_drive_out         : out   std_logic ;
    pwr_clock_out         : out   std_logic ;
    pwr_fpga_out          : out   std_logic ;
    pwr_sdram_out         : out   std_logic ;
    pwr_mram_out          : out   std_logic ;
    pwr_im_out            : out   std_logic ;
    pwr_gps_out           : out   std_logic ;
    pwr_datatx_out        : out   std_logic ;
    pwr_micR_out          : out   std_logic ;
    pwr_micL_out          : out   std_logic ;
    pwr_sdcard_out        : out   std_logic ;
    pwr_ls_1p8_out        : out   std_logic ;
    pwr_ls_3p3_out        : out   std_logic ;

    solar_max_in          : in    std_logic ;
    solar_on_in           : in    std_logic ;
    solar_run_out         : out   std_logic ;
	 
		gpio_1				    : out   std_logic ;
		gpio_2				    : out   std_logic ;
		gpio_3				    : out   std_logic ;
		gpio_4				    : out   std_logic ;
		gpio_5				    : out   std_logic ;
		gpio_6				    : out   std_logic ;
		gpio_7				    : out   std_logic ;
		gpio_8				    : out   std_logic ;

    forced_start_in       : in    std_logic ;
    fpga_fs_out           : out   std_logic ;
    rtc_alarm_in          : in    std_logic

  ) ;

end entity PowerController ;


architecture rtl of PowerController is

  --  FPGA state

  signal fpga_turnon              : std_logic := '0' ;
  signal fpga_activated           : std_logic := '0' ;
  signal fpga_powered             : std_logic := '0' ;
  signal fpga_running             : std_logic := '0' ;

  --  Status and Control Registers.

  signal statreg_changed          : std_logic ;
  signal PC_StatusReg             : std_logic_vector (StatusSignalsCnt_c-1
                                                      downto 0) ;
  signal PC_ControlReg            : std_logic_vector (ControlSignalsCnt_c-1
                                                      downto 0) ;
  signal PC_ControlSet            : std_logic ;
  signal PC_ControlUse            : std_logic := '0' ;

  signal pwr_fpga_shutdown        : std_logic ;

  --  SPI lines.

  signal spi_miso                 : std_logic ;

  --  Signals that are inverts of the input of tri-stated signals.

  signal spi_cs                   : std_logic ;
  signal fpga_fs                  : std_logic ;

  --  Parallel Flash Loader signals.

  signal pfl_flash_cs             : std_logic_vector (0 downto 0) ;
  signal pfl_flash_clk            : std_logic_vector (0 downto 0) ;
  signal pfl_data                 : std_logic_vector (0 downto 0) ;
  signal pfl_dclk                 : std_logic ;
  signal pfl_nconfig              : std_logic ;
  signal pfl_flash_req            : std_logic ;

  alias  pfl_flash_io0            : std_logic_vector (0 downto 0) is
                                    pfl_flash_data_io (0 downto 0) ;
  alias  pfl_flash_io1            : std_logic_vector (0 downto 0) is
                                    pfl_flash_data_io (1 downto 1) ;
  alias  pfl_flash_io2            : std_logic_vector (0 downto 0) is
                                    pfl_flash_data_io (2 downto 2) ;
  alias  pfl_flash_io3            : std_logic_vector (0 downto 0) is
                                    pfl_flash_data_io (3 downto 3) ;

  --  Parallel Flash Loader.

  component PFL is
    port
    (
      fpga_conf_done            : IN    STD_LOGIC ;
      fpga_nstatus              : IN    STD_LOGIC ;
      fpga_pgm                  : IN    STD_LOGIC_VECTOR (2 DOWNTO 0);
      pfl_clk                   : IN    STD_LOGIC ;
      pfl_flash_access_granted  : IN    STD_LOGIC ;
      pfl_nreset                : IN    STD_LOGIC ;
      flash_io0                 : INOUT STD_LOGIC_VECTOR (0 DOWNTO 0) ;
      flash_io1                 : INOUT STD_LOGIC_VECTOR (0 DOWNTO 0) ;
      flash_io2                 : INOUT STD_LOGIC_VECTOR (0 DOWNTO 0) ;
      flash_io3                 : INOUT STD_LOGIC_VECTOR (0 DOWNTO 0) ;
      flash_ncs                 : OUT   STD_LOGIC_VECTOR (0 DOWNTO 0) ;
      flash_sck                 : OUT   STD_LOGIC_VECTOR (0 DOWNTO 0) ;
      fpga_data                 : OUT   STD_LOGIC_VECTOR (0 DOWNTO 0) ;
      fpga_dclk                 : OUT   STD_LOGIC ;
      fpga_nconfig              : OUT   STD_LOGIC ;
      pfl_flash_access_request  : OUT   STD_LOGIC
    ) ;
  end component PFL ;

  --  Status/Control SPI to FPGA.

  component StatCtlSPI is

    Generic (
      status_bits_g           : natural := 1 ;
      control_bits_g          : natural := 1
    ) ;
    Port (
      clk                     : in    std_logic ;
      status_in               : in    std_logic_vector (status_bits_g-1
                                                        downto 0) ;
      status_chg_out          : out   std_logic ;
      control_out             : out   std_logic_vector (control_bits_g-1
                                                        downto 0) ;
      control_set_out         : out   std_logic ;
      enable_in               : in    std_logic ;
      data_in                 : in    std_logic ;
      data_out                : out   std_logic
    ) ;

  end component StatCtlSPI ;

begin

  --  When the FPGA is not running all outputs to it will be zero.
  --  When the FPGA is not powered all inputs from it will be driven zero.
  --  When it is powered they will be high impedence.
  --
  --  Thus, when the FPGA is powered down all lines going to it from the
  --  Power Controller will be 0V, preventing any current flow through
  --  the FPGA to them.
  --  When the FPGA is starting up it sets all its lines to high impedence
  --  with a weak pull-up resistor.  At his time the Power Controller sets
  --  all its input lines from the FPGA to high impedence without a weak
  --  pull-up.  This results in no current flow through these lines then
  --  and into the time the FPGA is running.

  master_clk_out        <= '0' when (fpga_running = '0') else master_clk ;

  flash_clk_out         <= pfl_flash_clk (0) when (fpga_running = '0') else
                           fpga_toflash_clk_in ;
  flash_cs_out          <= pfl_flash_cs  (0) when (fpga_running = '0') else
                           fpga_toflash_cs_in ;
  fpga_flash_data_io    <= "0000" when (fpga_powered = '0') else
                           "ZZZZ" when (fpga_running = '0') else
                           "ZZZZ" when (fpga_toflash_dir_in = '0') else
                           fpga_toflash_data_io ;
  fpga_toflash_data_io  <= "0000" when (fpga_powered = '0') else
                           "ZZZZ" when (fpga_running = '0') else
                           "ZZZZ" when (fpga_toflash_dir_in = '1') else
                           fpga_flash_data_io ;
  fpga_toflash_clk_in   <= '0' when (fpga_powered = '0') else 'Z' ;
  fpga_toflash_cs_in    <= '0' when (fpga_powered = '0') else 'Z' ;
  fpga_toflash_dir_in   <= '0' when (fpga_powered = '0') else 'Z' ;

  fpga_cnf_dclk_out     <= '0' when (fpga_powered = '0') else
                           pfl_dclk ;
  fpga_cnf_data_out     <= '0' when (fpga_powered = '0') else
                           pfl_data (0) ;
									
                  
                  
  --Debug--
  --This is the sequence of FPGA turn on events as conducted by the CPLD.
  gpio_1 					<=	fpga_activated;
  gpio_2 					<=	fpga_powered;
  gpio_3 					<=	fpga_running;
  --Debug--								

  fpga_cnf_nconfig_out  <= '1' when (fpga_activated = '0') else
                           pfl_nconfig ;

  statchg_out           <= '0' when (fpga_running = '0') else
                           statreg_changed ;
  spi_miso_out          <= '0' when (fpga_running = '0') else
                           spi_miso ;
  spi_clk_in            <= '0' when (fpga_powered = '0') else 'Z' ;
  spi_cs_in             <= '0' when (fpga_powered = '0') else 'Z' ;
  spi_cs                <= not spi_cs_in ;
  spi_mosi_in           <= '0' when (fpga_powered = '0') else 'Z' ;

  bat_int_fpga_out      <= '0' when (fpga_running = '0') else
                           bat_int_in ;
  fpga_fs_out           <= '0' when (fpga_running = '0') else
                           fpga_fs ;
  fpga_fs               <= not forced_start_in ;

  i2c_clk_io            <= 'Z' ;
  i2c_data_io           <= 'Z' ;

  --  Activate the Octal Buffer drive.

  pwr_drive_out         <= '1' ;

  --  Start the FPGA when a battery monitor interrupt occurs and the
  --  FPGA is not running.

  fpga_turnon           <= (not fpga_running) and
                           --(bat_int_in        or
                            --forced_start_in   or
                            --rtc_alarm_in
									 forced_start_in ;

  --  Devices powered as FPGA is starting.

  pwr_clock_out         <= '0' when (fpga_activated  = '0') else '1' ;

  pwr_pwm_out           <= '0' when (fpga_activated  = '0') else '1' ;

  pwr_2p5_run_out       <= '0' when (fpga_activated  = '0') else '1' ;
  pwr_3p3_run_out       <= '0' when (pwr_2p5_good_in = '0') else '1' ;
  pwr_1p1_run_out       <= '0' when (pwr_3p3_good_in = '0') else '1' ;

  pwr_fpga_out          <= '0' when (pwr_1p1_good_in = '0') else '1' ;

  fpga_running          <= '0' when (fpga_powered          = '0' or
                                     fpga_cnf_init_done_in = '0' or 
												  fpga_cnf_conf_done_in = '0' )
                               else '1' ;

  --  Status Register Bit Mappings.

  PC_StatusReg (StatusSignals'pos(Stat_BatteryGood_e))  <= bat_good_in ;
  PC_StatusReg (StatusSignals'pos(Stat_SolarCtlOn_e))   <= solar_on_in ;
  PC_StatusReg (StatusSignals'pos(Stat_SolarCtlMax_e))  <= solar_max_in ;
  PC_StatusReg (StatusSignals'pos(Stat_BattMonLow_e))   <= bat_low_in ;
  PC_StatusReg (StatusSignals'pos(Stat_ForceStartup_e)) <= forced_start_in ;
  PC_StatusReg (StatusSignals'pos(Stat_PwrGood2p5_e))   <= pwr_2p5_good_in ;
  PC_StatusReg (StatusSignals'pos(Stat_PwrGood3p3_e))   <= pwr_3p3_good_in ;
  PC_StatusReg (StatusSignals'pos(Stat_Spacer1_e))      <= '0' ;
  PC_StatusReg (StatusSignals'pos(Stat_Spacer2_e))      <= '0' ;

  --  Control Register Bit Mappings and default values.

  bat_power_out         <=
        PC_ControlReg (ControlSignals'pos(Ctl_MainPowerSwitch_e))
        when (PC_ControlUse = '1') else '1' ;
  bat_recharge_out      <=
        PC_ControlReg (ControlSignals'pos(Ctl_RechargeSwitch_e))
        when (PC_ControlUse = '1') else '1' ;
  solar_run_out         <=
        PC_ControlReg (ControlSignals'pos(Ctl_SolarCtlShutdown_e))
        when (PC_ControlUse = '1') else '0' ;
  pwr_ls_3p3_out        <=
        PC_ControlReg (ControlSignals'pos(Ctl_LevelShifter3p3_e))
        when (PC_ControlUse = '1') else '0' ;
  pwr_ls_1p8_out        <=
        PC_ControlReg (ControlSignals'pos(Ctl_LevelShifter1p8_e))
        when (PC_ControlUse = '1') else '0' ;
  pwr_im_out            <=
        PC_ControlReg (ControlSignals'pos(Ctl_InertialOn1p8_e))
        when (PC_ControlUse = '1') else '0' ;
  pwr_micL_out          <=
        PC_ControlReg (ControlSignals'pos(Ctl_MicLeftOn_e))
        when (PC_ControlUse = '1') else '0' ;
  pwr_micR_out          <=
        PC_ControlReg (ControlSignals'pos(Ctl_MicRightOn_e))
        when (PC_ControlUse = '1') else '0' ;
  pwr_sdram_out         <=
        PC_ControlReg (ControlSignals'pos(Ctl_SDRAM_On_e))
        when (PC_ControlUse = '1') else '0' ;
  pwr_sdcard_out        <=
        PC_ControlReg (ControlSignals'pos(Ctl_SDCardOn_e))
        when (PC_ControlUse = '1') else '0' ;
  pwr_mram_out          <=
        PC_ControlReg (ControlSignals'pos(Ctl_MagMemOn_e))
        when (PC_ControlUse = '1') else '0' ;
  pwr_gps_out           <=
        PC_ControlReg (ControlSignals'pos(Ctl_GPS_On_e))
        when (PC_ControlUse = '1') else '0' ;
  pwr_datatx_out        <=
        PC_ControlReg (ControlSignals'pos(Ctl_DataTX_On_e))
        when (PC_ControlUse = '1') else '0' ;
  pwr_fpga_shutdown     <=
        PC_ControlReg (ControlSignals'pos(Ctl_FPGA_Shutdown_e))
        when (PC_ControlUse = '1') else '0' ;

  --  Parallel Flash Loader.
  --  When pfl_flash_access_granted is low all flash_* lines are
  --  tri-stated.  (PFL Users Guide Table 15).  This prevents JTAG access
  --  to flash and FPGA configuration.  (PFL Users Guide Table 17).
  --  Hold the pfl_nreset low to prevent FPGA configuration.  (PFL Users
  --  Guide Table 15).  This does not prevent JTAG programming of flash.

  pfl_inst : PFL
    port map
    (
      fpga_conf_done            => fpga_cnf_conf_done_in,
      fpga_nstatus              => fpga_cnf_nstatus_in,
      fpga_pgm                  => "000",
      pfl_clk                   => master_clk,
      pfl_flash_access_granted  => '1',
      pfl_nreset                => (fpga_activated and not fpga_running),
      flash_io0                 => pfl_flash_io0,
      flash_io1                 => pfl_flash_io1,
      flash_io2                 => pfl_flash_io2,
      flash_io3                 => pfl_flash_io3,
      flash_ncs                 => pfl_flash_cs,
      flash_sck                 => pfl_flash_clk,
      fpga_data                 => pfl_data,
      fpga_dclk                 => pfl_dclk,
      fpga_nconfig              => pfl_nconfig,
      pfl_flash_access_request  => pfl_flash_req
    ) ;

  --  Status/Control SPI to FPGA.

  FPGA_SPI : StatCtlSPI

    Generic Map (
      status_bits_g           => PC_StatusReg'length,
      control_bits_g          => PC_ControlReg'length
    )
    Port Map (
      clk                     => not spi_clk_in,
      status_in               => PC_StatusReg,
      status_chg_out          => statreg_changed,
      control_out             => PC_ControlReg,
      control_set_out         => PC_ControlSet,
      enable_in               => not spi_cs,
      data_in                 => spi_mosi_in,
      data_out                => spi_miso
    ) ;

  --------------------------------------------------------------------------
  --  Turn the FPGA on and off based on the turnon and shutdown signals.
  --------------------------------------------------------------------------

  fpga_on_off : process (fpga_turnon, pwr_fpga_shutdown)
  begin
    if (fpga_turnon = '1') then
      fpga_activated    <= '1' ;

    elsif (rising_edge (pwr_fpga_shutdown)) then
      fpga_activated    <= '0' ;
    end if ;
  end process fpga_on_off ;


  --------------------------------------------------------------------------
  --  Set the FPGA powered condition when the FPGA responds that it is
  --  ready to be configured.
  --------------------------------------------------------------------------

  fpga_powerup : process (fpga_activated, fpga_cnf_nstatus_in)
  begin
    if (fpga_activated = '0') then
      fpga_powered      <= '0' ;

    elsif (rising_edge (fpga_cnf_nstatus_in)) then
      fpga_powered      <= '1' ;
    end if ;
  end process fpga_powerup ;


  --------------------------------------------------------------------------
  --  Set the control register value.
  --------------------------------------------------------------------------

  ctl_set : process (fpga_running, PC_ControlSet)
  begin
    if (fpga_running = '0') then
      PC_ControlUse     <= '0' ;

    elsif (rising_edge (PC_ControlSet)) then
      PC_ControlUse     <= '1' ;
    end if ;
  end process ctl_set ;


end architecture rtl ;
