-- megafunction wizard: %ALTUFM_NONE%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: ALTUFM_NONE 

-- ============================================================
-- File Name: Flash.vhd
-- Megafunction Name(s):
-- 			ALTUFM_NONE
--
-- Simulation Library Files(s):
-- 			maxv
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 13.1.0 Build 162 10/23/2013 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2013 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--altufm_none CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="MAX V" ERASE_TIME=500000000 OSC_FREQUENCY=180000 PORT_ARCLKENA="PORT_UNUSED" PORT_DRCLKENA="PORT_UNUSED" PROGRAM_TIME=1600000 WIDTH_UFM_ADDRESS=9 arclk ardin arshft busy drclk drdin drdout drshft erase osc oscena program rtpbusy
--VERSION_BEGIN 13.1 cbx_a_gray2bin 2013:10:23:18:05:48:SJ cbx_a_graycounter 2013:10:23:18:05:48:SJ cbx_altufm_none 2013:10:23:18:05:48:SJ cbx_cycloneii 2013:10:23:18:05:48:SJ cbx_lpm_add_sub 2013:10:23:18:05:48:SJ cbx_lpm_compare 2013:10:23:18:05:48:SJ cbx_lpm_counter 2013:10:23:18:05:48:SJ cbx_lpm_decode 2013:10:23:18:05:48:SJ cbx_lpm_mux 2013:10:23:18:05:48:SJ cbx_maxii 2013:10:23:18:05:48:SJ cbx_mgl 2013:10:23:18:06:54:SJ cbx_stratix 2013:10:23:18:05:48:SJ cbx_stratixii 2013:10:23:18:05:48:SJ cbx_util_mgl 2013:10:23:18:05:48:SJ  VERSION_END

 LIBRARY maxv;
 USE maxv.all;

--synthesis_resources = maxv_ufm 1 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  Flash_altufm_none_4bp IS 
	 PORT 
	 ( 
		 arclk	:	IN  STD_LOGIC;
		 ardin	:	IN  STD_LOGIC;
		 arshft	:	IN  STD_LOGIC;
		 busy	:	OUT  STD_LOGIC;
		 drclk	:	IN  STD_LOGIC;
		 drdin	:	IN  STD_LOGIC;
		 drdout	:	OUT  STD_LOGIC;
		 drshft	:	IN  STD_LOGIC;
		 erase	:	IN  STD_LOGIC;
		 osc	:	OUT  STD_LOGIC;
		 oscena	:	IN  STD_LOGIC;
		 program	:	IN  STD_LOGIC;
		 rtpbusy	:	OUT  STD_LOGIC
	 ); 
 END Flash_altufm_none_4bp;

 ARCHITECTURE RTL OF Flash_altufm_none_4bp IS

	 SIGNAL  wire_maxii_ufm_block1_bgpbusy	:	STD_LOGIC;
	 SIGNAL  wire_maxii_ufm_block1_busy	:	STD_LOGIC;
	 SIGNAL  wire_maxii_ufm_block1_drdout	:	STD_LOGIC;
	 SIGNAL  wire_maxii_ufm_block1_osc	:	STD_LOGIC;
	 SIGNAL  ufm_arclk :	STD_LOGIC;
	 SIGNAL  ufm_ardin :	STD_LOGIC;
	 SIGNAL  ufm_arshft :	STD_LOGIC;
	 SIGNAL  ufm_bgpbusy :	STD_LOGIC;
	 SIGNAL  ufm_busy :	STD_LOGIC;
	 SIGNAL  ufm_drclk :	STD_LOGIC;
	 SIGNAL  ufm_drdin :	STD_LOGIC;
	 SIGNAL  ufm_drdout :	STD_LOGIC;
	 SIGNAL  ufm_drshft :	STD_LOGIC;
	 SIGNAL  ufm_erase :	STD_LOGIC;
	 SIGNAL  ufm_osc :	STD_LOGIC;
	 SIGNAL  ufm_oscena :	STD_LOGIC;
	 SIGNAL  ufm_program :	STD_LOGIC;
	 COMPONENT  maxv_ufm
	 GENERIC 
	 (
		ADDRESS_WIDTH	:	NATURAL := 9;
		ERASE_TIME	:	NATURAL := 500000000;
		INIT_FILE	:	STRING := "UNUSED";
		mem1	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem10	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem11	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem12	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem13	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem14	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem15	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem16	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem2	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem3	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem4	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem5	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem6	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem7	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem8	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		mem9	:	STD_LOGIC_VECTOR(511 DOWNTO 0) := "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
		OSC_SIM_SETTING	:	NATURAL := 180000;
		PROGRAM_TIME	:	NATURAL := 1600000;
		lpm_type	:	STRING := "maxv_ufm"
	 );
	 PORT
	 ( 
		arclk	:	IN STD_LOGIC := '0';
		ardin	:	IN STD_LOGIC := '0';
		arshft	:	IN STD_LOGIC := '1';
		bgpbusy	:	OUT STD_LOGIC;
		busy	:	OUT STD_LOGIC;
		drclk	:	IN STD_LOGIC := '0';
		drdin	:	IN STD_LOGIC := '0';
		drdout	:	OUT STD_LOGIC;
		drshft	:	IN STD_LOGIC := '1';
		erase	:	IN STD_LOGIC := '0';
		osc	:	OUT STD_LOGIC;
		oscena	:	IN STD_LOGIC := '0';
		program	:	IN STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
 BEGIN

	busy <= ufm_busy;
	drdout <= ufm_drdout;
	osc <= ufm_osc;
	rtpbusy <= ufm_bgpbusy;
	ufm_arclk <= arclk;
	ufm_ardin <= ardin;
	ufm_arshft <= arshft;
	ufm_bgpbusy <= wire_maxii_ufm_block1_bgpbusy;
	ufm_busy <= wire_maxii_ufm_block1_busy;
	ufm_drclk <= drclk;
	ufm_drdin <= drdin;
	ufm_drdout <= wire_maxii_ufm_block1_drdout;
	ufm_drshft <= drshft;
	ufm_erase <= erase;
	ufm_osc <= wire_maxii_ufm_block1_osc;
	ufm_oscena <= oscena;
	ufm_program <= program;
	maxii_ufm_block1 :  maxv_ufm
	  GENERIC MAP (
		ADDRESS_WIDTH => 9,
		ERASE_TIME => 500000000,
		INIT_FILE => "none",
		mem1 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem10 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem11 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem12 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem13 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem14 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem15 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem16 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem2 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem3 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem4 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem5 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem6 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem7 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem8 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		mem9 => "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
		OSC_SIM_SETTING => 180000,
		PROGRAM_TIME => 1600000
	  )
	  PORT MAP ( 
		arclk => ufm_arclk,
		ardin => ufm_ardin,
		arshft => ufm_arshft,
		bgpbusy => wire_maxii_ufm_block1_bgpbusy,
		busy => wire_maxii_ufm_block1_busy,
		drclk => ufm_drclk,
		drdin => ufm_drdin,
		drdout => wire_maxii_ufm_block1_drdout,
		drshft => ufm_drshft,
		erase => ufm_erase,
		osc => wire_maxii_ufm_block1_osc,
		oscena => ufm_oscena,
		program => ufm_program
	  );

 END RTL; --Flash_altufm_none_4bp
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY Flash IS
	PORT
	(
		arclk		: IN STD_LOGIC ;
		ardin		: IN STD_LOGIC ;
		arshft		: IN STD_LOGIC ;
		drclk		: IN STD_LOGIC ;
		drdin		: IN STD_LOGIC ;
		drshft		: IN STD_LOGIC ;
		erase		: IN STD_LOGIC ;
		oscena		: IN STD_LOGIC ;
		program		: IN STD_LOGIC ;
		busy		: OUT STD_LOGIC ;
		drdout		: OUT STD_LOGIC ;
		osc		: OUT STD_LOGIC ;
		rtpbusy		: OUT STD_LOGIC 
	);
END Flash;


ARCHITECTURE RTL OF flash IS

	SIGNAL sub_wire0	: STD_LOGIC ;
	SIGNAL sub_wire1	: STD_LOGIC ;
	SIGNAL sub_wire2	: STD_LOGIC ;
	SIGNAL sub_wire3	: STD_LOGIC ;



	COMPONENT Flash_altufm_none_4bp
	PORT (
			arshft	: IN STD_LOGIC ;
			drclk	: IN STD_LOGIC ;
			erase	: IN STD_LOGIC ;
			program	: IN STD_LOGIC ;
			arclk	: IN STD_LOGIC ;
			drdin	: IN STD_LOGIC ;
			osc	: OUT STD_LOGIC ;
			oscena	: IN STD_LOGIC ;
			rtpbusy	: OUT STD_LOGIC ;
			ardin	: IN STD_LOGIC ;
			drdout	: OUT STD_LOGIC ;
			busy	: OUT STD_LOGIC ;
			drshft	: IN STD_LOGIC 
	);
	END COMPONENT;

BEGIN
	osc    <= sub_wire0;
	rtpbusy    <= sub_wire1;
	drdout    <= sub_wire2;
	busy    <= sub_wire3;

	Flash_altufm_none_4bp_component : Flash_altufm_none_4bp
	PORT MAP (
		arshft => arshft,
		drclk => drclk,
		erase => erase,
		program => program,
		arclk => arclk,
		drdin => drdin,
		oscena => oscena,
		ardin => ardin,
		drshft => drshft,
		osc => sub_wire0,
		rtpbusy => sub_wire1,
		drdout => sub_wire2,
		busy => sub_wire3
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "MAX V"
-- Retrieval info: CONSTANT: ERASE_TIME NUMERIC "500000000"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "MAX V"
-- Retrieval info: CONSTANT: LPM_FILE STRING "UNUSED"
-- Retrieval info: CONSTANT: LPM_HINT STRING "UNUSED"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altufm_none"
-- Retrieval info: CONSTANT: OSC_FREQUENCY NUMERIC "180000"
-- Retrieval info: CONSTANT: PORT_ARCLKENA STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_DRCLKENA STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PROGRAM_TIME NUMERIC "1600000"
-- Retrieval info: CONSTANT: WIDTH_UFM_ADDRESS NUMERIC "9"
-- Retrieval info: USED_PORT: arclk 0 0 0 0 INPUT NODEFVAL "arclk"
-- Retrieval info: CONNECT: @arclk 0 0 0 0 arclk 0 0 0 0
-- Retrieval info: USED_PORT: ardin 0 0 0 0 INPUT NODEFVAL "ardin"
-- Retrieval info: CONNECT: @ardin 0 0 0 0 ardin 0 0 0 0
-- Retrieval info: USED_PORT: arshft 0 0 0 0 INPUT NODEFVAL "arshft"
-- Retrieval info: CONNECT: @arshft 0 0 0 0 arshft 0 0 0 0
-- Retrieval info: USED_PORT: busy 0 0 0 0 OUTPUT NODEFVAL "busy"
-- Retrieval info: CONNECT: busy 0 0 0 0 @busy 0 0 0 0
-- Retrieval info: USED_PORT: drclk 0 0 0 0 INPUT NODEFVAL "drclk"
-- Retrieval info: CONNECT: @drclk 0 0 0 0 drclk 0 0 0 0
-- Retrieval info: USED_PORT: drdin 0 0 0 0 INPUT NODEFVAL "drdin"
-- Retrieval info: CONNECT: @drdin 0 0 0 0 drdin 0 0 0 0
-- Retrieval info: USED_PORT: drdout 0 0 0 0 OUTPUT NODEFVAL "drdout"
-- Retrieval info: CONNECT: drdout 0 0 0 0 @drdout 0 0 0 0
-- Retrieval info: USED_PORT: drshft 0 0 0 0 INPUT NODEFVAL "drshft"
-- Retrieval info: CONNECT: @drshft 0 0 0 0 drshft 0 0 0 0
-- Retrieval info: USED_PORT: erase 0 0 0 0 INPUT NODEFVAL "erase"
-- Retrieval info: CONNECT: @erase 0 0 0 0 erase 0 0 0 0
-- Retrieval info: USED_PORT: osc 0 0 0 0 OUTPUT NODEFVAL "osc"
-- Retrieval info: CONNECT: osc 0 0 0 0 @osc 0 0 0 0
-- Retrieval info: USED_PORT: oscena 0 0 0 0 INPUT NODEFVAL "oscena"
-- Retrieval info: CONNECT: @oscena 0 0 0 0 oscena 0 0 0 0
-- Retrieval info: USED_PORT: program 0 0 0 0 INPUT NODEFVAL "program"
-- Retrieval info: CONNECT: @program 0 0 0 0 program 0 0 0 0
-- Retrieval info: USED_PORT: rtpbusy 0 0 0 0 OUTPUT NODEFVAL "rtpbusy"
-- Retrieval info: CONNECT: rtpbusy 0 0 0 0 @rtpbusy 0 0 0 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL Flash.vhd TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Flash.qip TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Flash.bsf FALSE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Flash_inst.vhd FALSE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Flash.inc FALSE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Flash.cmp FALSE TRUE
-- Retrieval info: LIB_FILE: maxv
