----------------------------------------------------------------------------
--
--! @file       Collar.vhd
--! @brief      Acoustic Recording Collar Top Level.
--! @details    Instanciates and connects all the components that make up the
--!             Acoustic Recording Collar FPGA implementation.
--! @author     Emery Newlon
--! @date       August 2014
--! @copyright  Copyright (C) 2014 Ross K. Snider and Emery L. Newlon
--
--  This program is free software: you can redistribute it and/or modify
--  it under the terms of the GNU General Public License as published by
--  the Free Software Foundation, either version 3 of the License, or
--  (at your option) any later version.
--
--  This program is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--  GNU General Public License for more details.
--
--  You should have received a copy of the GNU General Public License
--  along with this program.  If not, see <http://www.gnu.org/licenses/>.
--
--  Emery Newlon
--  Electrical and Computer Engineering
--  Montana State University
--  610 Cobleigh Hall
--  Bozeman, MT 59717
--  emery.newlon@msu.montana.edu
--
----------------------------------------------------------------------------

library IEEE ;                  --! Use standard library.
use IEEE.STD_LOGIC_1164.ALL ;   --! Use standard logic elements.
use IEEE.NUMERIC_STD.ALL ;      --! Use numeric standard.
use IEEE.MATH_REAL.ALL ;        --! Real number functions.

library GENERAL ;               --! General libraries
use GENERAL.UTILITIES_PKG.ALL ;

use GENERAL.GPS_CLOCK_PKG.ALL ;

library WORK ;                  --! Local Library
use WORK.COLLAR_CONTROL_PKG.ALL ;


----------------------------------------------------------------------------
--
--! @brief      Acoustic Recording Collar Top Level.
--! @details    Instanciates and connects all the components that make up
--!             the Acoustic Recording Collar FPGA implementation.
--!
--! @param      master_clk_freq_g Frequency of the system clock in cycles
--!                               per second.
--! @param      button_cnt_g    Number of buttons used by the device.
--! @param      master_clk      Clock generated by the system that drives
--!                             everything else.
--! @param      buttons_in      Vector of button signals used by the device.
--! @param      batt_int_in     Battery monitor interrupt signal.
--! @param      forced_start_in A forced startup has been initiated.
--! @param      i2c_clk_io      I2C bus clock is input or output depending
--!                             on the device driving it.
--! @param      i2c_data_io     I2C bus data is driven by the same device
--!                             that is driving the clock.
--! @param      pc_statchg_in   The Power Controller status register has
--!                             changed and should be reloaded.
--! @param      pc_spi_clk      The Power Controller status register/
--!                             control register SPI bus clock.
--! @param      pc_spi_cs_out   The PC SPI bus chip select.  An SPI
--!                             transfer is initiated when it goes high.
--! @param      pc_spi_mosi_out Master Out/Slave In SPI data line.
--! @param      pc_spi_miso_in  Master In/Slave Out SPI data line.
--! @param      pc_flash_clk      Power Controller Flash access clock.
--! @param      pc_flash_cs_out   PC Flash chip select.
--! @param      pc_flash_data_io  PC Flash data bus.
--! @param      pc_flash_dir_out  PC Flash data direction.  The PC Flash
--!                               bus is high impedance when this line is
--!                               low, driven when it is high.
--! @param      sdram_clk         Clock driving the SDRAM.
--! @param      sdram_clk_en_out  The clock is enabled on the SDRAM.
--! @param      sdram_command_out The command sent to the SDRAM.
--! @param      sdram_mask_out    The bytes masked from the SDRAM data bus.
--! @param      sdram_bank_out    The SDRAM bank to access.
--! @param      sdram_addr_out    The SDRAM row or column to access.
--! @param      sdram_data_io     The SDRAM data bus.
--! @param      sd_clk          Micro SDCard clock.
--! @param      sd_cmd_io       Command line used with the micro SDCard.
--! @param      sd_data_io      Data lines used with the micro SDCard.
--! @param      sd_vsw_out      Voltage switch control lines.
--! @param      sdh_clk         High voltage micro SDCard clock.
--! @param      sdh_cmd_io      High voltage command line used with the
--!                             micro SDCard.
--! @param      sdh_data_io     High voltage data lines used with the micro
--!                             SDCard.
--! @param      gps_rx_in       Receive line from the GPS UART.
--! @param      gps_tx_out      Transmit line to the GPS UART.
--! @param      gps_timemark_out  Time mark generator line to the GPS external
--!                               interrupt.
--! @param      ms_clk          Motion sensor SPI Clock.
--! @param      ms_cs_out       Motion sensor SPI chip select.
--! @param      ms_mosi_out     Motion sensor SPI Master Out/Slave In.
--! @param      ms_miso_in      Motion sensor SPI Master In/Slave Out.
--! @param      ms_int_in       Motion sensor Interrupt.
--! @param      ms_cs_accgyro_out   Motion sensor A/G SPI chip select.
--! @param      ms_miso_accgyro_in  Motion sensor A/G SPI Master In/Slave
--!                                 Out.
--! @param      ms_int1_accgyro_in  Motion sensor A/G Interrupt 1.
--! @param      ms_int2_accgyro_in  Motion sensor A/G Interrupt 2.
--! @param      ms_cs_mag_out   Motion sensor magnetic SPI chip select.
--! @param      ms_miso_mag_in  Motion sensor magnetic SPI Master In/
--!                             Slave Out.
--! @param      ms_int_mag_in   Motion sensor magnetic Interrupt.
--! @param      ms_drdy_mag_in  Motion sensor magnetic Data Ready.
--! @param      magram_clk            Magnetic RAM SPI clock.
--! @param      magram_cs_out         Magnetic RAM chip select.
--! @param      magram_mosi_out       Magnetic RAM SPI Master Out/Slave In.
--! @param      magram_miso_in        Magnetic RAM SPI Master In/Slave Out.
--! @param      magram_writeprot_out  Magnetic RAM write protect.
--! @param      mic_clk         Microphone clock.
--! @param      mic_right_in    Right microphone data.
--! @param      mic_left_in     Left microphone data.
--! @param      radio_clk       Radio trx/rcv bus clock.
--! @param      radio_data_io   Radio data bus.
--
----------------------------------------------------------------------------

entity Collar is

  Generic (
    master_clk_freq_g     : natural   := 10e6 ;
    button_cnt_g          : natural   :=  8
  ) ;
  Port (
    master_clk            : in    std_logic ;
    buttons_in            : in    std_logic_vector (button_cnt_g-1
                                                      downto 0) ;

    batt_int_in           : in    std_logic ;
    forced_start_in       : in    std_logic ;

    i2c_clk_io            : inout std_logic ;
    i2c_data_io           : inout std_logic ;

    pc_statchg_in         : in    std_logic ;
    pc_spi_clk            : out   std_logic ;
    pc_spi_cs_out         : out   std_logic ;
    pc_spi_mosi_out       : out   std_logic ;
    pc_spi_miso_in        : in    std_logic ;

    pc_flash_clk          : out   std_logic ;
    pc_flash_cs_out       : out   std_logic ;
    pc_flash_data_io      : inout std_logic_vector (3 downto 0) ;
    pc_flash_dir_out      : out   std_logic ;

    sdram_clk             : out   std_logic ;
    sdram_clk_en_out      : out   std_logic ;
    sdram_command_out     : out   std_logic_vector (3 downto 0) ;
    sdram_mask_out        : out   std_logic_vector (1 downto 0) ;
    sdram_bank_out        : out   std_logic_vector (1 downto 0) ;
    sdram_addr_out        : out   std_logic_vector (13 downto 0) ;
    sdram_data_io         : inout std_logic_vector (15 downto 0) ;

    sd_clk                : out   std_logic ;
    sd_cmd_io             : inout std_logic ;
    sd_data_io            : inout std_logic_vector (3 downto 0) ;
    sd_vsw_out            : out   std_logic_vector (1 downto 0) ;

    sdh_clk               : out   std_logic ;
    sdh_cmd_io            : inout std_logic ;
    sdh_data_io           : inout std_logic_vector (3 downto 0) ;

    gps_rx_in             : in    std_logic ;
    gps_tx_out            : out   std_logic ;
    gps_timemark_out      : out   std_logic ;

    ms_clk                : out   std_logic ;
    ms_cs_out             : out   std_logic ;
    ms_mosi_out           : out   std_logic ;
    ms_miso_in            : in    std_logic ;
    ms_int_in             : in    std_logic ;

    ms_cs_accgyro_out     : out   std_logic ;
    ms_miso_accgyro_in    : in    std_logic ;
    ms_int1_accgyro_in    : in    std_logic ;
    ms_int2_accgyro_in    : in    std_logic ;

    ms_cs_mag_out         : out   std_logic ;
    ms_miso_mag_in        : in    std_logic ;
    ms_int_mag_in         : in    std_logic ;
    ms_drdy_mag_in        : in    std_logic ;

    magram_clk            : out   std_logic ;
    magram_cs_out         : out   std_logic ;
    magram_mosi_out       : out   std_logic ;
    magram_miso_in        : in    std_logic ;
    magram_writeprot_out  : out   std_logic ;

    mic_clk               : out   std_logic ;
    mic_right_in          : in    std_logic ;
    mic_left_in           : in    std_logic ;

    radio_clk             : out   std_logic ;
    radio_data_io         : inout std_logic_vector (4 downto 0)
  ) ;

end entity Collar ;


architecture structural of Collar is

  --  Button specifications.

  constant reset_button_c     : natural := 0 ;
  constant sd_start_button_c  : natural := 1 ;

  --  Reset clock signals.

  signal reset_time         : GPS_Time ;

  --  Reset information.  The power up signal defaults to zero.

  constant pb_time_c        : real    := 0.5 ;
  constant pb_count_c       : natural :=
              natural (trunc (real (master_clk_freq_g) * pb_time_c)) ;
  constant pb_count_bits_c  : natural := const_bits (pb_count_c) ;

  signal reset              : std_logic ;
  signal power_up           : std_logic := '0' ;
  signal reset_pushed       : std_logic := '0' ;
  signal pb_counter         : unsigned (pb_count_bits_c-1 downto 0) :=
                                (others => '0') ;

  --  GPS signals.

  signal aop_running        : std_logic ;

  --  GPS dual port RAM communication signals.

  constant gpsmemsrc_addrbits_c : natural := 9 ;
  constant gpsmemsrc_databits_c : natural := 8 ;

  signal gpsmemsrc_addr         : std_logic_vector (gpsmemsrc_addrbits_c-1
                                                    downto 0) ;
  signal gpsmemsrc_clk          : std_logic ;
  signal gpsmemsrc_writeto      : std_logic_vector (gpsmemsrc_databits_c-1
                                                    downto 0) ;
  signal gpsmemsrc_readfrom     : std_logic_vector (gpsmemsrc_databits_c-1
                                                    downto 0) ;
  signal gpsmemsrc_read_en      : std_logic ;
  signal gpsmemsrc_write_en     : std_logic ;

  constant gpsmemdst_addrbits_c : natural := 9 ;
  constant gpsmemdst_databits_c : natural := 8 ;

  signal gpsmemdst_addr         : std_logic_vector (gpsmemdst_addrbits_c-1
                                                    downto 0) ;
  signal gpsmemdst_clk          : std_logic ;
  signal gpsmemdst_readfrom     : std_logic_vector (gpsmemdst_databits_c-1
                                                    downto 0) ;
  signal gpsmemdst_read_en      : std_logic ;
  signal gpsmemdst_write_en     : std_logic ;

  constant gps_baudrate_c       : natural := 9600 ;

  --  Clock specifications.

  constant gps_clk_freq_c     : natural := gps_baudrate_c * 16 ;
  constant gps_clk_cntmax_c   : natural := master_clk_freq_g /
                                           (gps_clk_freq_c * 2) ;

  constant gps_clk_cntbits_c  : natural := const_bits (gps_clk_cntmax_c) ;

  signal gps_clk_cnt          : unsigned (gps_clk_cntbits_c-1 downto 0) ;

  signal gps_clk              : std_logic ;

begin

  --------------------------------------------------------------------------
  --  Time since reset clock.
  --------------------------------------------------------------------------

  use_StrClk:
    if (Collar_Control_useStrClk_c = '1') generate

      component StartupClock is

        Generic (
          CLK_FREQ              : natural := 50e6
        ) ;
        Port (
          clk                   : in    std_logic ;
          time_since_reset_out  : out   GPS_Time
        ) ;

      end component StartupClock ;

    begin

      reset_clock : StartupClock
        Generic Map (
          CLK_FREQ              => master_clk_freq_g
        )
        Port Map (
          clk                   => master_clk,
          time_since_reset_out  => reset_time
        ) ;

  end generate use_StrClk ;

  --------------------------------------------------------------------------
  --  I2C bus.
  --------------------------------------------------------------------------

  no_use_I2C:
    if (Collar_Control_useI2C_c = '0') generate

      i2c_clk_io              <= '0' ;
      i2c_data_io             <= '0' ;

    end generate no_use_I2c ;

  --------------------------------------------------------------------------
  --  Power Controller.
  --------------------------------------------------------------------------

  no_use_PC:
    if (Collar_Control_usePC_c = '0') generate

      pc_spi_clk              <= '0' ;
      pc_spi_cs_out           <= '1' ;
      pc_spi_mosi_out         <= '0' ;

      pc_flash_clk            <= '0' ;
      pc_flash_cs_out         <= '1' ;
      pc_flash_data_io        <= (others => 'Z') ;
      pc_flash_dir_out        <= '0' ;

    end generate no_use_PC ;

  --------------------------------------------------------------------------
  --  SDRAM.
  --------------------------------------------------------------------------

  no_use_SDRAM:
    if (Collar_Control_useSDRAM_c = '0') generate

      sdram_clk               <= '0' ;
      sdram_clk_en_out        <= '0' ;
      sdram_command_out       <= (others => '1') ;
      sdram_mask_out          <= (others => '0') ;
      sdram_bank_out          <= (others => '0') ;
      sdram_addr_out          <= (others => '0') ;
      sdram_data_io           <= (others => '0') ;

    end generate no_use_SDRAM ;

  --------------------------------------------------------------------------
  --  SD Card controller.
  --------------------------------------------------------------------------

  use_SD:
    if (Collar_Control_useSD_c = '1') generate

      component microsd_controller is
        generic (
          BUFSIZE         : natural   := 2048 ;
          HS_SDR25_MODE   : std_logic := '1' ;
          CLK_DIVIDE      : natural   := 128
        ) ;
        port (
          rst_n           : in    std_logic ;
          clk             : in    std_logic ;
          clock_enable    : in    std_logic ;

          data_input      : in    std_logic_vector (7 downto 0) ;
          data_we         : in    std_logic ;
          data_full       : out   std_logic ;

          data_sd_start_address : in    std_logic_vector (31 downto 0) ;
          data_nblocks          : in    std_logic_vector (31 downto 0) ;

          sd_clk          : out   std_logic ;
          sd_cmd          : inout std_logic ;
          sd_dat          : inout std_logic_vector (3 downto 0) ;

          V_3_3_ON_OFF    : out   std_logic ;
          V_1_8_ON_OFF    : out   std_logic ;

          init_start      : in    std_logic ;
          user_led_n_out  : out   std_logic_vector (3 downto 0)
        ) ;
      end component microsd_controller ;

    begin

      sdcard : microsd_controller
        generic map (
          BUFSIZE         => 2048,
          HS_SDR25_MODE   => '1',
          CLK_DIVIDE      => natural (real (master_clk_freq_g) / 400000.0)
        )
        port map (
          rst_n           => not reset,
          clk             => master_clk,
          clock_enable    => '0',

          data_input      => (others => '0'),
          data_we         => '0',

          data_sd_start_address => (others => '0'),
          data_nblocks          => (others => '0'),

          sd_clk          => sd_clk,
          sd_cmd          => sd_cmd_io,
          sd_dat          => sd_data_io,

          V_3_3_ON_OFF    => sd_vsw_out (0),
          V_1_8_ON_OFF    => sd_vsw_out (1),

          init_start      => '0'
        ) ;

    end generate use_SD ;

  no_use_SD:
    if (Collar_Control_useSD_c = '0') generate

      sd_clk        <= '0' ;
      sd_cmd_io     <= '0' ;
      sd_data_io    <= (others => '0') ;
      sd_vsw_out    <= (others => '0') ;

    end generate no_use_SD ;

  --------------------------------------------------------------------------
  --  Direct connect SD Card controller.  Does not use voltage level
  --  shifting.
  --------------------------------------------------------------------------

  use_SDH:
    if (Collar_Control_useSDH_c = '1') generate

      component microsd_controller is
        generic (
          BUFSIZE         : natural   := 2048 ;
          HS_SDR25_MODE   : std_logic := '1' ;
          CLK_DIVIDE      : natural   := 128
        ) ;
        port (
          rst_n           : in    std_logic ;
          clk             : in    std_logic ;
          clock_enable    : in    std_logic ;

          data_input      : in    std_logic_vector (7 downto 0) ;
          data_we         : in    std_logic ;
          data_full       : out   std_logic ;

          data_sd_start_address : in    std_logic_vector (31 downto 0) ;
          data_nblocks          : in    std_logic_vector (31 downto 0) ;

          sd_clk          : out   std_logic ;
          sd_cmd          : inout std_logic ;
          sd_dat          : inout std_logic_vector (3 downto 0) ;

          V_3_3_ON_OFF    : out   std_logic ;
          V_1_8_ON_OFF    : out   std_logic ;

          init_start      : in    std_logic ;
          user_led_n_out  : out   std_logic_vector (3 downto 0)
        ) ;
      end component microsd_controller ;

    begin

      sdcard : microsd_controller
        generic map (
          BUFSIZE         => 2048,
          HS_SDR25_MODE   => '1',
          CLK_DIVIDE      => natural (real (master_clk_freq_g) / 400000.0)
        )
        port map (
          rst_n           => not reset,
          clk             => master_clk,
          clock_enable    => '0',

          data_input      => (others => '0'),
          data_we         => '0',

          data_sd_start_address => (others => '0'),
          data_nblocks          => (others => '0'),

          sd_clk          => sdh_clk,
          sd_cmd          => sdh_cmd_io,
          sd_dat          => sdh_data_io,

          init_start      => '0'
        ) ;

  end generate use_SDH ;

  no_use_SDH:
    if (Collar_Control_useSDH_c = '0') generate

      sdh_clk        <= '0' ;
      sdh_cmd_io     <= '0' ;
      sdh_data_io    <= (others => '0') ;

  end generate no_use_SDH ;

  --------------------------------------------------------------------------
  --  GPS RAM
  --------------------------------------------------------------------------

  use_GPS_RAM:
    if (Collar_Control_useGPS_c = '1') generate

      component gps_ram IS
        PORT
        (
          address_a		: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
          address_b		: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
          clock_a		: IN STD_LOGIC  := '1';
          clock_b		: IN STD_LOGIC ;
          data_a		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
          data_b		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
          rden_a		: IN STD_LOGIC  := '1';
          rden_b		: IN STD_LOGIC  := '1';
          wren_a		: IN STD_LOGIC  := '0';
          wren_b		: IN STD_LOGIC  := '0';
          q_a		: OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
          q_b		: OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
        );
      END component gps_ram;

    begin

      --  Memory component.  Clock is triggered on negative going edge to allow
      --  input signals to propagate in one half clock cycle and to produce
      --  output by the next clock cycle.  The memory is fast enough to produce
      --  output in less than one half clock cycle.

      gps_ramblocks : gps_ram
        Port Map (
          address_a		            => gpsmemsrc_addr,
          address_b		            => gpsmemdst_addr,
          clock_a		              => gpsmemsrc_clk,
          clock_b		              => gpsmemdst_clk,
          data_a		              => gpsmemsrc_writeto,
          data_b		              => (others => '0'),
          rden_a		              => gpsmemsrc_read_en,
          rden_b		              => gpsmemdst_read_en,
          wren_a		              => gpsmemsrc_write_en,
          wren_b		              => '0',
          q_a		                  => gpsmemsrc_readfrom,
          q_b		                  => gpsmemdst_readfrom
        ) ;

  end generate use_GPS_RAM ;

  no_use_GPS_RAM:
    if (Collar_Control_useGPS_c = '0') generate

      gpsmemsrc_addr      <= (others => '0') ;
      gpsmemsrc_clk       <= '0' ;
      gpsmemsrc_writeto   <= (others => '0') ;
      gpsmemsrc_read_en   <= '0' ;
      gpsmemsrc_write_en  <= '0' ;

      gpsmemdst_addr      <= (others => '0') ;
      gpsmemdst_clk       <= '0' ;
      gpsmemdst_read_en   <= '0' ;

  end generate no_use_GPS_RAM ;

  --------------------------------------------------------------------------
  --  GPS Message controller.
  --------------------------------------------------------------------------

  use_GPS:
    if (Collar_Control_useGPS_c = '1') generate

      component GPSmessages is

        Generic (
          clk_freq_g            : natural := 50e6 ;
          mem_addrbits_g        : natural := 9 ;
          mem_databits_g        : natural := 8
        ) ;
        Port (
          reset                 : in    std_logic ;
          clk                   : in    std_logic ;
          curtime_in            : in    std_logic_vector (gps_time_bits_c-1
                                                          downto 0) ;
          pollinterval_in       : in    unsigned (13 downto 0) ;
          gpsmem_clk_out        : out   std_logic ;
          gpsmem_addr_out       : out   std_logic_vector (mem_addrbits_g-1
                                                          downto 0) ;
          gpsmem_read_en_out    : out   std_logic ;
          gpsmem_write_en_out   : out   std_logic ;
          gpsmem_readfrom_in    : in    std_logic_vector (mem_databits_g-1
                                                          downto 0) ;
          gpsmem_writeto_out    : out   std_logic_vector (mem_databits_g-1
                                                          downto 0) ;
          gps_rx_in             : in    std_logic ;
          gps_tx_out            : out   std_logic ;
          timemarker_out        : out   std_logic ;
          aop_running_out       : out   std_logic
        ) ;

      end component GPSmessages ;

      --  GPS control signals.

      signal poll_int         : unsigned (13 downto 0) :=
                                        TO_UNSIGNED (15, 14) ;

    begin

      gps_ctl : GPSmessages
        Generic Map (
          clk_freq_g            => gps_clk_freq_c,
          mem_addrbits_g        => gpsmemsrc_addrbits_c,
          mem_databits_g        => gpsmemsrc_databits_c
        )
        Port (
          reset                 => reset,
          clk                   => gps_clk,
          curtime_in            => reset_time,
          pollinterval_in       => poll_int,
          gpsmem_clk_out        => gpsmemsrc_clk,
          gpsmem_addr_out       => gpsmemsrc_addr,
          gpsmem_read_en_out    => gpsmemsrc_read_en,
          gpsmem_write_en_out   => gpsmemsrc_write_en,
          gpsmem_readfrom_in    => gpsmemsrc_readfrom,
          gpsmem_writeto_out    => gpsmemsrc_writeto,
          gps_rx                => gps_rx_in,
          gps_tx                => gps_tx_out,
          timemarker            => gps_timemark_out,
          aop_running_out       => aop_running
        ) ;

  end generate use_GPS ;

  no_use_GPS:
    if (Collar_Control_useGPS_c = '0') generate

      gps_tx_out        <= '0' ;
      gps_timemark_out  <= '0' ;
      aop_running       <= '0' ;

  end generate no_use_GPS ;

  --------------------------------------------------------------------------
  --  Inertial sensor controller.
  --------------------------------------------------------------------------

  no_use_Inertial:
    if (Collar_Control_useInertial_c = '0') generate

      ms_clk                  <= '0' ;
      ms_cs_out               <= '1' ;
      ms_mosi_out             <= '0' ;

      ms_cs_accgyro_out       <= '1' ;

      ms_cs_mag_out           <= '1' ;

    end generate no_use_Inertial ;

  --------------------------------------------------------------------------
  --  Magnetic RAM control.
  --------------------------------------------------------------------------

  no_use_MagMem:
    if (Collar_Control_useMagMem_c = '0') generate

      magram_clk              <= '0' ;
      magram_cs_out           <= '1' ;
      magram_mosi_out         <= '0' ;
      magram_writeprot_out    <= '0' ;

    end generate no_use_MagMem ;

  --------------------------------------------------------------------------
  --  Microphone control.
  --------------------------------------------------------------------------

  no_use_PDMmic:
    if (Collar_Control_usePDMmic_c = '0') generate

      mic_clk                 <= '0' ;

    end generate no_use_PDMmic ;

  --------------------------------------------------------------------------
  --  Radio control.
  --------------------------------------------------------------------------

  no_use_Radio:
    if (Collar_Control_useRadio_c = '0') generate

      radio_clk               <= '0' ;
      radio_data_io           <= (others => '0') ;

    end generate no_use_Radio ;


  --------------------------------------------------------------------------
  --  Reset occurs on power up or button press of the reset button.
  --------------------------------------------------------------------------

  reset                     <= (not power_up) or reset_pushed ;

  reset_poweron : process (master_clk)
  begin
    if (rising_edge (master_clk)) then
      power_up              <= '1' ;
    end if ;
  end process reset_poweron ;

  --  Debounce the reset button by making sure it is held up or down for a
  --  long period of time.

  reset_pb : process (master_clk)
  begin
    if (rising_edge (master_clk)) then

      if (buttons_in (reset_button_c) /= reset_pushed) then
        if (pb_counter = pb_count_c) then
          reset_pushed      <= buttons_in (reset_button_c) ;
          pb_counter        <= (others => '0') ;
        else
          pb_counter        <= pb_counter + 1 ;
        end if ;
      else
        pb_counter          <= (others => '0') ;
      end if ;
    end if ;
  end process reset_pb ;

  --------------------------------------------------------------------------
  --  GPS clock generation.
  --------------------------------------------------------------------------

  gps_clk_gen : process (reset, master_clk)
  begin
    if (reset = '1') then
      gps_clk_cnt     <= (others => '0') ;
      gps_clk         <= '0' ;

    elsif (rising_edge (master_clk)) then
      if (gps_clk_cnt /= TO_UNSIGNED (gps_clk_cntmax_c,
                                      gps_clk_cnt'length)) then

        gps_clk_cnt  <= gps_clk_cnt + 1 ;
      else
        gps_clk_cnt  <= (others => '0') ;
        gps_clk      <= not gps_clk;
      end if ;
    end if ;

  end process gps_clk_gen ;

end architecture structural ;
