----------------------------------------------------------------------------
--
--! @file       PowerController.vhd
--! @brief      Power Controller Top Level.
--! @details    Instanciates and connects all the components that make up
--!             the Power Controller CPLD implementation.
--! @author     Emery Newlon
--! @date       September 2014
--! @copyright  Copyright (C) 2014 Ross K. Snider and Emery L. Newlon
--
--  This program is free software: you can redistribute it and/or modify
--  it under the terms of the GNU General Public License as published by
--  the Free Software Foundation, either version 3 of the License, or
--  (at your option) any later version.
--
--  This program is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--  GNU General Public License for more details.
--
--  You should have received a copy of the GNU General Public License
--  along with this program.  If not, see <http://www.gnu.org/licenses/>.
--
--  Emery Newlon
--  Electrical and Computer Engineering
--  Montana State University
--  610 Cobleigh Hall
--  Bozeman, MT 59717
--  emery.newlon@msu.montana.edu
--
----------------------------------------------------------------------------

library IEEE ;                  --! Use standard library.
use IEEE.STD_LOGIC_1164.ALL ;   --! Use standard logic elements.
use IEEE.NUMERIC_STD.ALL ;      --! Use numeric standard.
use IEEE.MATH_REAL.ALL ;        --! Real number functions.

library GENERAL ;               --! General libraries
use GENERAL.UTILITIES_PKG.ALL ;


----------------------------------------------------------------------------
--
--! @brief      Power Controller Top Level.
--! @details    Instanciates and connects all the components that make up
--!             the Power Controller CPLD implementation.
--!
--! @param      master_clk_freq_g Frequency of the system clock in cycles
--!                               per second.
--! @param      master_clk        Clock generated by the system that drives
--!                               everything else.
--! @param      master_clk_out    Output of the master clock to the FPGA.
--!
--! @param      flash_clk_out         Flash clock.
--! @param      flash_cs_out          Flash chip select.
--! @param      pfl_flash_data_io     Parallel Flash Loader Flash data bus.
--! @param      fpga_flash_data_io    FPGA Flash data bus.
--! @param      fpga_toflash_clk_in   FPGA to Flash clock.
--! @param      fpga_toflash_cs_in    FPGA to Flash chip select.
--! @param      fpga_toflash_data_io  FPGA to Flash data bus.
--! @param      fpga_toflash_dir_in   FPGA to Flash data direction.
--!
--! @param      fpga_cnf_dclk_out     FPGA Configuration data clock.
--! @param      fpga_cnf_data_out     FPGA Configuration data to FPGA.
--! @param      fpga_cnf_nstatus_in   FPGA Configuration status not.
--! @param      fpga_cnf_conf_done_in FPGA Configuration config done.
--! @param      fpga_cnf_init_done_in FPGA Configuration init done.
--! @param      fpga_cnf_nconfig_out  FPGA Configuration configure not.
--!
--! @param      statchg_out       The status register has changed.
--! @param      spi_clk_in        The PC status register / FPGA control
--!                               register SPI bus clock.
--! @param      spi_cs_in         The PC SPI bus chip select.  An SPI
--!                               transfer is initiated when it goes high.
--! @param      spi_mosi_in       Master Out/Slave In SPI data line.
--! @param      spi_miso_out      Master In/Slave Out SPI data line.
--!
--! @param      i2c_clk_io        I2C bus clock is input or output depending
--!                               on the device driving it.
--! @param      i2c_data_io       I2C bus data is driven by the same device
--!                               that is driving the clock.
--!
--! @param      bat_power_out     Battery power switch.
--! @param      bat_recharge_out  Battery recharge switch.
--! @param      bat_int_in        Battery monitor interrupt.
--! @param      bat_int_fpga_out  Battery monitor interrupt to FPGA.
--! @param      bat_low_in        Battery monitor battery low.
--! @param      bat_good_in       Battery monitor battery good.
--!
--! @param      pwr_1p1_run_out   Power on the 1.1 V power supply.
--! @param      pwr_1p1_good_in   The 1.1 V power supply is operating.
--! @param      pwr_2p5_run_out   Power on the 2.5 V power supply.
--! @param      pwr_2p5_good_in   The 2.5 V power supply is operating.
--! @param      pwr_3p3_run_out   Power on the 3.3 V power supply.
--! @param      pwr_3p3_good_in   The 3.3 V power supply is operating.
--! @param      pwr_pwm_out       Use PWM or burst mode.
--!
--! @param      pwr_drive_out     Drive the power switch buffer signals.
--! @param      pwr_clock_out     Power on the clock.
--! @param      pwr_fpga_out      Power on the FPGA 1.8, 2.5, & 3.3 Vcc.
--! @param      pwr_sdram_out     Power on the SDRAM.
--! @param      pwr_mram_out      Power on the Magnetic RAM.
--! @param      pwr_im_out        Power on the Inertial Modules.
--! @param      pwr_gps_out       Power on the GPS.
--! @param      pwr_datatx_out    Power on the Data Transmitter.
--! @param      pwr_micR_out      Power on the Right Hand Microphone.
--! @param      pwr_micL_out      Power on the Left Hand Microphone.
--! @param      pwr_sdcard_out    Power on the SD Cards.
--! @param      pwr_ls_1p8_out    Power on the 1.8 V Level Shifter.
--! @param      pwr_ls_3p3_out    Power on the 3.3 V Level Shifter.
--!
--! @param      solar_max_in      Solar Controller voltage level is at max.
--! @param      solar_on_in       Solar Controller is operating.
--! @param      solar_run_out     Solar Controller is turned on.
--!
--! @param      forced_start_in   A forced startup has been initiated.
--! @param      fpga_fs_out       Forced startup passed to the FPGA.
--! @param      rtc_alarm_in      Alarm interrupt from the Real Time Clock.
--
----------------------------------------------------------------------------

entity PowerController is

  Generic (
    master_clk_freq_g     : natural   := 10e6
  ) ;
  Port (
    master_clk            : in    std_logic ;
    master_clk_out        : out   std_logic ;

    flash_clk_out         : out   std_logic ;
    flash_cs_out          : out   std_logic ;
    pfl_flash_data_io     : inout std_logic_vector (3 downto 0) ;
    fpga_flash_data_io    : inout std_logic_vector (3 downto 0) ;
    fpga_toflash_clk_in   : in    std_logic ;
    fpga_toflash_cs_in    : in    std_logic ;
    fpga_toflash_data_io  : inout std_logic_vector (3 downto 0) ;
    fpga_toflash_dir_in   : in    std_logic ;

    fpga_cnf_dclk_out     : out   std_logic ;
    fpga_cnf_data_out     : out   std_logic ;
    fpga_cnf_nstatus_in   : in    std_logic ;
    fpga_cnf_conf_done_in : in    std_logic ;
    fpga_cnf_init_done_in : in    std_logic ;
    fpga_cnf_nconfig_out  : out   std_logic ;

    statchg_out           : out   std_logic ;
    spi_clk_in            : in    std_logic ;
    spi_cs_in             : in    std_logic ;
    spi_mosi_in           : in    std_logic ;
    spi_miso_out          : out   std_logic ;

    i2c_clk_io            : inout std_logic ;
    i2c_data_io           : inout std_logic ;

    bat_power_out         : out   std_logic ;
    bat_recharge_out      : out   std_logic ;
    bat_int_in            : in    std_logic ;
    bat_int_fpga_out      : out   std_logic ;
    bat_low_in            : in    std_logic ;
    bat_good_in           : in    std_logic ;

    pwr_1p1_run_out       : out   std_logic ;
    pwr_1p1_good_in       : in    std_logic ;
    pwr_2p5_run_out       : out   std_logic ;
    pwr_2p5_good_in       : in    std_logic ;
    pwr_3p3_run_out       : out   std_logic ;
    pwr_3p3_good_in       : in    std_logic ;
    pwr_pwm_out           : out   std_logic ;

    pwr_drive_out         : out   std_logic ;
    pwr_clock_out         : out   std_logic ;
    pwr_fpga_out          : out   std_logic ;
    pwr_sdram_out         : out   std_logic ;
    pwr_mram_out          : out   std_logic ;
    pwr_im_out            : out   std_logic ;
    pwr_gps_out           : out   std_logic ;
    pwr_datatx_out        : out   std_logic ;
    pwr_micR_out          : out   std_logic ;
    pwr_micL_out          : out   std_logic ;
    pwr_sdcard_out        : out   std_logic ;
    pwr_ls_1p8_out        : out   std_logic ;
    pwr_ls_3p3_out        : out   std_logic ;

    solar_max_in          : in    std_logic ;
    solar_on_in           : in    std_logic ;
    solar_run_out         : out   std_logic ;

    forced_start_in       : in    std_logic ;
    fpga_fs_out           : out   std_logic ;
    rtc_alarm_in          : in    std_logic

  ) ;

end entity PowerController ;


architecture structural of PowerController is

  --  FPGA state

  signal fpga_running             : std_logic := '0' ;


begin

  --  When the FPGA is not running all outputs to it will be zero.  All
  --  inputs from it will be high impedence.

  master_clk_out        <= '0' when (fpga_running = '0') else master_clk ;

  flash_clk_out         <= pfl_flash_clk when (fpga_running = '0') else
                           fpga_toflash_clk_in ;
  flash_cs_out          <= pfl_flash_cs  when (fpga_running = '0') else
                           fpga_toflash_cs_in ;
  fpga_flash_data_io    <= 'Z' when (fpga_running = '0') else
                           'Z' when (fpga_toflash_dir_in = '0') else
                           fpga_toflash_data_io ;
  fpga_toflash_data_io  <= '0' when (fpga_running = '0') else
                           'Z' when (fpga_toflash_dir_in = '1') else
                           fpga_flash_data_io ;

  fpga_cnf_dclk_out     <= '0' when (fpga_running = '0') else
                           pfl_dclk ;
  fpga_cnf_data_out     <= '0' when (fpga_running = '0') else
                           pfl_data ;
  fpga_cnf_nconfig_out  <= '0' when (fpga_running = '0') else
                           pfl_nconfig ;

  statchg_out           <= '0' when (fpga_running = '0') else
                           statreg_changed ;
  spi_miso_out          <= '0' when (fpga_running = '0') else
                           spi_miso ;

  bat_int_fpga_out      <= '0' when (fpga_running = '0') else
                           bat_int_in ;
  fpga_fs_out           <= '0' when (fpga_running = '0') else
                           forced_start_in ;


end architecture structural ;
